<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-2.16385,-13.2909,56.5218,-42.8443</PageViewport>
<gate>
<ID>2</ID>
<type>AA_LABEL</type>
<position>28.5,-11.5</position>
<gparam>LABEL_TEXT 1-bit register</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3</ID>
<type>AA_LABEL</type>
<position>7.5,-37.5</position>
<gparam>LABEL_TEXT Combinational Logic</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>AA_MUX_2x1</type>
<position>12,-25</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>1 </output>
<input>
<ID>SEL_0</ID>2 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_LABEL</type>
<position>30,-37.5</position>
<gparam>LABEL_TEXT Sequential Logic</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AE_DFF_LOW</type>
<position>30,-24</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>12 </output>
<input>
<ID>clock</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>10,-19</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>4,-24</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>20</ID>
<type>BB_CLOCK</type>
<position>23,-33</position>
<output>
<ID>CLK</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>22</ID>
<type>GA_LED</type>
<position>47,-22</position>
<input>
<ID>N_in0</ID>12 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>AA_LABEL</type>
<position>10,-16</position>
<gparam>LABEL_TEXT load</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>AA_LABEL</type>
<position>30.5,-18.5</position>
<gparam>LABEL_TEXT data-flip-flop</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>AA_LABEL</type>
<position>4,-21.5</position>
<gparam>LABEL_TEXT in</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>AA_LABEL</type>
<position>47,-25</position>
<gparam>LABEL_TEXT out</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24,-22,27,-22</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>24 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>24,-25,24,-22</points>
<intersection>-25 5</intersection>
<intersection>-22 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>14,-25,24,-25</points>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<intersection>24 4</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12,-22.5,12,-19</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<connection>
<GID>4</GID>
<name>SEL_0</name></connection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>6,-24,10,-24</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27,-33,27,-25</points>
<connection>
<GID>20</GID>
<name>CLK</name></connection>
<connection>
<GID>10</GID>
<name>clock</name></connection></vsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>10,-29.5,36,-29.5</points>
<intersection>10 5</intersection>
<intersection>36 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>36,-29.5,36,-22</points>
<intersection>-29.5 1</intersection>
<intersection>-22 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>33,-22,46,-22</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<connection>
<GID>22</GID>
<name>N_in0</name></connection>
<intersection>36 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>10,-29.5,10,-26</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>-29.5 1</intersection></vsegment></shape></wire></page 0>
<page 1>
<PageViewport>-139.611,2.09853,447.246,-293.435</PageViewport>
<gate>
<ID>33</ID>
<type>AA_LABEL</type>
<position>34.5,-7</position>
<gparam>LABEL_TEXT 16-bits register</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>AA_MUX_2x1</type>
<position>35.5,-23.5</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>15 </input>
<output>
<ID>OUT</ID>13 </output>
<input>
<ID>SEL_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>35</ID>
<type>AE_DFF_LOW</type>
<position>46.5,-25.5</position>
<input>
<ID>IN_0</ID>13 </input>
<output>
<ID>OUT_0</ID>17 </output>
<input>
<ID>clock</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_TOGGLE</type>
<position>16,-17.5</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>37</ID>
<type>AA_TOGGLE</type>
<position>27.5,-22.5</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>38</ID>
<type>BB_CLOCK</type>
<position>-3,-147</position>
<output>
<ID>CLK</ID>69 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>39</ID>
<type>GA_LED</type>
<position>58,-23.5</position>
<input>
<ID>N_in0</ID>17 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>AA_LABEL</type>
<position>15.5,-14.5</position>
<gparam>LABEL_TEXT load</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>41</ID>
<type>AA_LABEL</type>
<position>46.5,-19.5</position>
<gparam>LABEL_TEXT data-flip-flop</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>AA_LABEL</type>
<position>27.5,-20</position>
<gparam>LABEL_TEXT in[0]</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>43</ID>
<type>AA_LABEL</type>
<position>58,-25.5</position>
<gparam>LABEL_TEXT out[0]</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>50</ID>
<type>AA_MUX_2x1</type>
<position>35,-38.5</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>22 </input>
<output>
<ID>OUT</ID>21 </output>
<input>
<ID>SEL_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>51</ID>
<type>AE_DFF_LOW</type>
<position>46,-40.5</position>
<input>
<ID>IN_0</ID>21 </input>
<output>
<ID>OUT_0</ID>23 </output>
<input>
<ID>clock</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>52</ID>
<type>AA_TOGGLE</type>
<position>27,-37.5</position>
<output>
<ID>OUT_0</ID>22 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>53</ID>
<type>GA_LED</type>
<position>57.5,-38.5</position>
<input>
<ID>N_in0</ID>23 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>54</ID>
<type>AA_LABEL</type>
<position>27,-35</position>
<gparam>LABEL_TEXT in[1]</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>55</ID>
<type>AA_LABEL</type>
<position>57.5,-40.5</position>
<gparam>LABEL_TEXT out[1]</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>56</ID>
<type>AA_MUX_2x1</type>
<position>34.5,-53</position>
<input>
<ID>IN_0</ID>26 </input>
<input>
<ID>IN_1</ID>25 </input>
<output>
<ID>OUT</ID>24 </output>
<input>
<ID>SEL_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>57</ID>
<type>AE_DFF_LOW</type>
<position>45.5,-55</position>
<input>
<ID>IN_0</ID>24 </input>
<output>
<ID>OUT_0</ID>26 </output>
<input>
<ID>clock</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>58</ID>
<type>AA_TOGGLE</type>
<position>26.5,-52</position>
<output>
<ID>OUT_0</ID>25 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>59</ID>
<type>GA_LED</type>
<position>57,-53</position>
<input>
<ID>N_in0</ID>26 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>AA_LABEL</type>
<position>26.5,-49.5</position>
<gparam>LABEL_TEXT in[2]</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>61</ID>
<type>AA_LABEL</type>
<position>57,-55</position>
<gparam>LABEL_TEXT out[2]</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>62</ID>
<type>AA_MUX_2x1</type>
<position>34.5,-69</position>
<input>
<ID>IN_0</ID>29 </input>
<input>
<ID>IN_1</ID>28 </input>
<output>
<ID>OUT</ID>27 </output>
<input>
<ID>SEL_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>63</ID>
<type>AE_DFF_LOW</type>
<position>45.5,-71</position>
<input>
<ID>IN_0</ID>27 </input>
<output>
<ID>OUT_0</ID>29 </output>
<input>
<ID>clock</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>64</ID>
<type>AA_TOGGLE</type>
<position>26.5,-68</position>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>65</ID>
<type>GA_LED</type>
<position>57,-69</position>
<input>
<ID>N_in0</ID>29 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>66</ID>
<type>AA_LABEL</type>
<position>26.5,-65.5</position>
<gparam>LABEL_TEXT in[3]</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>67</ID>
<type>AA_LABEL</type>
<position>57,-71</position>
<gparam>LABEL_TEXT out[3]</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>68</ID>
<type>AA_MUX_2x1</type>
<position>34,-84</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>31 </input>
<output>
<ID>OUT</ID>30 </output>
<input>
<ID>SEL_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>69</ID>
<type>AE_DFF_LOW</type>
<position>45,-86</position>
<input>
<ID>IN_0</ID>30 </input>
<output>
<ID>OUT_0</ID>32 </output>
<input>
<ID>clock</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>70</ID>
<type>AA_TOGGLE</type>
<position>26,-83</position>
<output>
<ID>OUT_0</ID>31 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>71</ID>
<type>GA_LED</type>
<position>56.5,-84</position>
<input>
<ID>N_in0</ID>32 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>72</ID>
<type>AA_LABEL</type>
<position>26,-80.5</position>
<gparam>LABEL_TEXT in[3]</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>73</ID>
<type>AA_LABEL</type>
<position>56.5,-86</position>
<gparam>LABEL_TEXT out[3]</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>74</ID>
<type>AA_MUX_2x1</type>
<position>33.5,-98.5</position>
<input>
<ID>IN_0</ID>35 </input>
<input>
<ID>IN_1</ID>34 </input>
<output>
<ID>OUT</ID>33 </output>
<input>
<ID>SEL_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>75</ID>
<type>AE_DFF_LOW</type>
<position>44.5,-100.5</position>
<input>
<ID>IN_0</ID>33 </input>
<output>
<ID>OUT_0</ID>35 </output>
<input>
<ID>clock</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>76</ID>
<type>AA_TOGGLE</type>
<position>25.5,-97.5</position>
<output>
<ID>OUT_0</ID>34 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>77</ID>
<type>GA_LED</type>
<position>56,-98.5</position>
<input>
<ID>N_in0</ID>35 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>78</ID>
<type>AA_LABEL</type>
<position>25.5,-95</position>
<gparam>LABEL_TEXT in[4]</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>79</ID>
<type>AA_LABEL</type>
<position>56,-100.5</position>
<gparam>LABEL_TEXT out[4]</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>80</ID>
<type>AA_MUX_2x1</type>
<position>33,-111.5</position>
<input>
<ID>IN_0</ID>38 </input>
<input>
<ID>IN_1</ID>37 </input>
<output>
<ID>OUT</ID>36 </output>
<input>
<ID>SEL_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>81</ID>
<type>AE_DFF_LOW</type>
<position>44,-113.5</position>
<input>
<ID>IN_0</ID>36 </input>
<output>
<ID>OUT_0</ID>38 </output>
<input>
<ID>clock</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>82</ID>
<type>AA_TOGGLE</type>
<position>25,-110.5</position>
<output>
<ID>OUT_0</ID>37 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>83</ID>
<type>GA_LED</type>
<position>55.5,-111.5</position>
<input>
<ID>N_in0</ID>38 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>84</ID>
<type>AA_LABEL</type>
<position>25,-108</position>
<gparam>LABEL_TEXT in[5]</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>85</ID>
<type>AA_LABEL</type>
<position>55.5,-113.5</position>
<gparam>LABEL_TEXT out[5]</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>86</ID>
<type>AA_MUX_2x1</type>
<position>33,-125.5</position>
<input>
<ID>IN_0</ID>41 </input>
<input>
<ID>IN_1</ID>40 </input>
<output>
<ID>OUT</ID>39 </output>
<input>
<ID>SEL_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>87</ID>
<type>AE_DFF_LOW</type>
<position>44,-127.5</position>
<input>
<ID>IN_0</ID>39 </input>
<output>
<ID>OUT_0</ID>41 </output>
<input>
<ID>clock</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>88</ID>
<type>AA_TOGGLE</type>
<position>25,-124.5</position>
<output>
<ID>OUT_0</ID>40 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>89</ID>
<type>GA_LED</type>
<position>55.5,-125.5</position>
<input>
<ID>N_in0</ID>41 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>90</ID>
<type>AA_LABEL</type>
<position>25,-122</position>
<gparam>LABEL_TEXT in[6]</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>91</ID>
<type>AA_LABEL</type>
<position>55.5,-127.5</position>
<gparam>LABEL_TEXT out[6]</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>92</ID>
<type>AA_MUX_2x1</type>
<position>32.5,-139.5</position>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>IN_1</ID>43 </input>
<output>
<ID>OUT</ID>42 </output>
<input>
<ID>SEL_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>93</ID>
<type>AE_DFF_LOW</type>
<position>43.5,-141.5</position>
<input>
<ID>IN_0</ID>42 </input>
<output>
<ID>OUT_0</ID>44 </output>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>94</ID>
<type>AA_TOGGLE</type>
<position>24.5,-138.5</position>
<output>
<ID>OUT_0</ID>43 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>95</ID>
<type>GA_LED</type>
<position>55,-139.5</position>
<input>
<ID>N_in0</ID>44 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>96</ID>
<type>AA_LABEL</type>
<position>24.5,-136</position>
<gparam>LABEL_TEXT in[7]</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>97</ID>
<type>AA_LABEL</type>
<position>55,-141.5</position>
<gparam>LABEL_TEXT out[7]</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>98</ID>
<type>AA_MUX_2x1</type>
<position>32.5,-153</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>46 </input>
<output>
<ID>OUT</ID>45 </output>
<input>
<ID>SEL_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>99</ID>
<type>AE_DFF_LOW</type>
<position>43.5,-155</position>
<input>
<ID>IN_0</ID>45 </input>
<output>
<ID>OUT_0</ID>47 </output>
<input>
<ID>clock</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>100</ID>
<type>AA_TOGGLE</type>
<position>24.5,-152</position>
<output>
<ID>OUT_0</ID>46 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>101</ID>
<type>GA_LED</type>
<position>55,-153</position>
<input>
<ID>N_in0</ID>47 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>102</ID>
<type>AA_LABEL</type>
<position>24.5,-149.5</position>
<gparam>LABEL_TEXT in[8]</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>103</ID>
<type>AA_LABEL</type>
<position>55,-155</position>
<gparam>LABEL_TEXT out[8]</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>104</ID>
<type>AA_MUX_2x1</type>
<position>33,-169</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>49 </input>
<output>
<ID>OUT</ID>48 </output>
<input>
<ID>SEL_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>105</ID>
<type>AE_DFF_LOW</type>
<position>44,-171</position>
<input>
<ID>IN_0</ID>48 </input>
<output>
<ID>OUT_0</ID>50 </output>
<input>
<ID>clock</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>106</ID>
<type>AA_TOGGLE</type>
<position>25,-168</position>
<output>
<ID>OUT_0</ID>49 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>107</ID>
<type>GA_LED</type>
<position>55.5,-169</position>
<input>
<ID>N_in0</ID>50 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>108</ID>
<type>AA_LABEL</type>
<position>25,-165.5</position>
<gparam>LABEL_TEXT in[9]</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>109</ID>
<type>AA_LABEL</type>
<position>55.5,-171</position>
<gparam>LABEL_TEXT out[9]</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>110</ID>
<type>AA_MUX_2x1</type>
<position>32.5,-183.5</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>52 </input>
<output>
<ID>OUT</ID>51 </output>
<input>
<ID>SEL_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>111</ID>
<type>AE_DFF_LOW</type>
<position>43.5,-185.5</position>
<input>
<ID>IN_0</ID>51 </input>
<output>
<ID>OUT_0</ID>53 </output>
<input>
<ID>clock</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>112</ID>
<type>AA_TOGGLE</type>
<position>24.5,-182.5</position>
<output>
<ID>OUT_0</ID>52 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>113</ID>
<type>GA_LED</type>
<position>55,-183.5</position>
<input>
<ID>N_in0</ID>53 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>114</ID>
<type>AA_LABEL</type>
<position>24.5,-180</position>
<gparam>LABEL_TEXT in[10]</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>115</ID>
<type>AA_LABEL</type>
<position>55,-185.5</position>
<gparam>LABEL_TEXT out[10]</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>116</ID>
<type>AA_MUX_2x1</type>
<position>32.5,-199.5</position>
<input>
<ID>IN_0</ID>56 </input>
<input>
<ID>IN_1</ID>55 </input>
<output>
<ID>OUT</ID>54 </output>
<input>
<ID>SEL_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>117</ID>
<type>AE_DFF_LOW</type>
<position>43.5,-201.5</position>
<input>
<ID>IN_0</ID>54 </input>
<output>
<ID>OUT_0</ID>56 </output>
<input>
<ID>clock</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>118</ID>
<type>AA_TOGGLE</type>
<position>24.5,-198.5</position>
<output>
<ID>OUT_0</ID>55 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>119</ID>
<type>GA_LED</type>
<position>55,-199.5</position>
<input>
<ID>N_in0</ID>56 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>120</ID>
<type>AA_LABEL</type>
<position>24.5,-196</position>
<gparam>LABEL_TEXT in[11]</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>121</ID>
<type>AA_LABEL</type>
<position>55,-201.5</position>
<gparam>LABEL_TEXT out[11]</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>122</ID>
<type>AA_MUX_2x1</type>
<position>30.5,-215.5</position>
<input>
<ID>IN_0</ID>59 </input>
<input>
<ID>IN_1</ID>58 </input>
<output>
<ID>OUT</ID>57 </output>
<input>
<ID>SEL_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>123</ID>
<type>AE_DFF_LOW</type>
<position>41.5,-217.5</position>
<input>
<ID>IN_0</ID>57 </input>
<output>
<ID>OUT_0</ID>59 </output>
<input>
<ID>clock</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>124</ID>
<type>AA_TOGGLE</type>
<position>22.5,-214.5</position>
<output>
<ID>OUT_0</ID>58 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>125</ID>
<type>GA_LED</type>
<position>53,-215.5</position>
<input>
<ID>N_in0</ID>59 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>126</ID>
<type>AA_LABEL</type>
<position>22.5,-212</position>
<gparam>LABEL_TEXT in[12]</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>127</ID>
<type>AA_LABEL</type>
<position>53,-217.5</position>
<gparam>LABEL_TEXT out[12]</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>128</ID>
<type>AA_MUX_2x1</type>
<position>32,-232</position>
<input>
<ID>IN_0</ID>62 </input>
<input>
<ID>IN_1</ID>61 </input>
<output>
<ID>OUT</ID>60 </output>
<input>
<ID>SEL_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>129</ID>
<type>AE_DFF_LOW</type>
<position>43,-234</position>
<input>
<ID>IN_0</ID>60 </input>
<output>
<ID>OUT_0</ID>62 </output>
<input>
<ID>clock</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>130</ID>
<type>AA_TOGGLE</type>
<position>24,-231</position>
<output>
<ID>OUT_0</ID>61 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>131</ID>
<type>GA_LED</type>
<position>54.5,-232</position>
<input>
<ID>N_in0</ID>62 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>132</ID>
<type>AA_LABEL</type>
<position>24,-228.5</position>
<gparam>LABEL_TEXT in[13]</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>133</ID>
<type>AA_LABEL</type>
<position>54.5,-234</position>
<gparam>LABEL_TEXT out[13]</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>134</ID>
<type>AA_MUX_2x1</type>
<position>31,-248</position>
<input>
<ID>IN_0</ID>65 </input>
<input>
<ID>IN_1</ID>64 </input>
<output>
<ID>OUT</ID>63 </output>
<input>
<ID>SEL_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>135</ID>
<type>AE_DFF_LOW</type>
<position>42,-250</position>
<input>
<ID>IN_0</ID>63 </input>
<output>
<ID>OUT_0</ID>65 </output>
<input>
<ID>clock</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>136</ID>
<type>AA_TOGGLE</type>
<position>23,-247</position>
<output>
<ID>OUT_0</ID>64 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>137</ID>
<type>GA_LED</type>
<position>53.5,-248</position>
<input>
<ID>N_in0</ID>65 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>138</ID>
<type>AA_LABEL</type>
<position>23,-244.5</position>
<gparam>LABEL_TEXT in[14]</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>139</ID>
<type>AA_LABEL</type>
<position>53.5,-250</position>
<gparam>LABEL_TEXT out[14]</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>140</ID>
<type>AA_MUX_2x1</type>
<position>32,-263</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>67 </input>
<output>
<ID>OUT</ID>66 </output>
<input>
<ID>SEL_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>141</ID>
<type>AE_DFF_LOW</type>
<position>43,-265</position>
<input>
<ID>IN_0</ID>66 </input>
<output>
<ID>OUT_0</ID>68 </output>
<input>
<ID>clock</ID>69 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>142</ID>
<type>AA_TOGGLE</type>
<position>24,-262</position>
<output>
<ID>OUT_0</ID>67 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>143</ID>
<type>GA_LED</type>
<position>54.5,-263</position>
<input>
<ID>N_in0</ID>68 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>144</ID>
<type>AA_LABEL</type>
<position>24,-259.5</position>
<gparam>LABEL_TEXT in[15]</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>145</ID>
<type>AA_LABEL</type>
<position>54.5,-265</position>
<gparam>LABEL_TEXT out[15]</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37.5,-23.5,43.5,-23.5</points>
<connection>
<GID>34</GID>
<name>OUT</name></connection>
<connection>
<GID>35</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>18,-257.5,18,-17.5</points>
<intersection>-257.5 33</intersection>
<intersection>-243 34</intersection>
<intersection>-227 31</intersection>
<intersection>-210 28</intersection>
<intersection>-194 30</intersection>
<intersection>-178.5 25</intersection>
<intersection>-163.5 23</intersection>
<intersection>-148.5 26</intersection>
<intersection>-134.5 19</intersection>
<intersection>-121 20</intersection>
<intersection>-107 21</intersection>
<intersection>-93.5 16</intersection>
<intersection>-79 11</intersection>
<intersection>-64.5 14</intersection>
<intersection>-48.5 15</intersection>
<intersection>-33.5 7</intersection>
<intersection>-17.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>18,-17.5,35.5,-17.5</points>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection>
<intersection>18 0</intersection>
<intersection>35.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>35.5,-21,35.5,-17.5</points>
<connection>
<GID>34</GID>
<name>SEL_0</name></connection>
<intersection>-17.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>18,-33.5,35,-33.5</points>
<intersection>18 0</intersection>
<intersection>35 9</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>35,-36,35,-33.5</points>
<connection>
<GID>50</GID>
<name>SEL_0</name></connection>
<intersection>-33.5 7</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>18,-79,34,-79</points>
<intersection>18 0</intersection>
<intersection>34 47</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>18,-64.5,34.5,-64.5</points>
<intersection>18 0</intersection>
<intersection>34.5 48</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>18,-48.5,34.5,-48.5</points>
<intersection>18 0</intersection>
<intersection>34.5 49</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>18,-93.5,33.5,-93.5</points>
<intersection>18 0</intersection>
<intersection>33.5 46</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>18,-134.5,32.5,-134.5</points>
<intersection>18 0</intersection>
<intersection>32.5 43</intersection></hsegment>
<hsegment>
<ID>20</ID>
<points>18,-121,33,-121</points>
<intersection>18 0</intersection>
<intersection>33 44</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>18,-107,33,-107</points>
<intersection>18 0</intersection>
<intersection>33 45</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>18,-163.5,33,-163.5</points>
<intersection>18 0</intersection>
<intersection>33 41</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>18,-178.5,32.5,-178.5</points>
<intersection>18 0</intersection>
<intersection>32.5 40</intersection></hsegment>
<hsegment>
<ID>26</ID>
<points>18,-148.5,32.5,-148.5</points>
<intersection>18 0</intersection>
<intersection>32.5 42</intersection></hsegment>
<hsegment>
<ID>28</ID>
<points>18,-210,30.5,-210</points>
<intersection>18 0</intersection>
<intersection>30.5 38</intersection></hsegment>
<hsegment>
<ID>30</ID>
<points>18,-194,32.5,-194</points>
<intersection>18 0</intersection>
<intersection>32.5 39</intersection></hsegment>
<hsegment>
<ID>31</ID>
<points>18,-227,32,-227</points>
<intersection>18 0</intersection>
<intersection>32 37</intersection></hsegment>
<hsegment>
<ID>33</ID>
<points>18,-257.5,32,-257.5</points>
<intersection>18 0</intersection>
<intersection>32 35</intersection></hsegment>
<hsegment>
<ID>34</ID>
<points>18,-243,31,-243</points>
<intersection>18 0</intersection>
<intersection>31 36</intersection></hsegment>
<vsegment>
<ID>35</ID>
<points>32,-260.5,32,-257.5</points>
<connection>
<GID>140</GID>
<name>SEL_0</name></connection>
<intersection>-257.5 33</intersection></vsegment>
<vsegment>
<ID>36</ID>
<points>31,-245.5,31,-243</points>
<connection>
<GID>134</GID>
<name>SEL_0</name></connection>
<intersection>-243 34</intersection></vsegment>
<vsegment>
<ID>37</ID>
<points>32,-229.5,32,-227</points>
<connection>
<GID>128</GID>
<name>SEL_0</name></connection>
<intersection>-227 31</intersection></vsegment>
<vsegment>
<ID>38</ID>
<points>30.5,-213,30.5,-210</points>
<connection>
<GID>122</GID>
<name>SEL_0</name></connection>
<intersection>-210 28</intersection></vsegment>
<vsegment>
<ID>39</ID>
<points>32.5,-197,32.5,-194</points>
<connection>
<GID>116</GID>
<name>SEL_0</name></connection>
<intersection>-194 30</intersection></vsegment>
<vsegment>
<ID>40</ID>
<points>32.5,-181,32.5,-178.5</points>
<connection>
<GID>110</GID>
<name>SEL_0</name></connection>
<intersection>-178.5 25</intersection></vsegment>
<vsegment>
<ID>41</ID>
<points>33,-166.5,33,-163.5</points>
<connection>
<GID>104</GID>
<name>SEL_0</name></connection>
<intersection>-163.5 23</intersection></vsegment>
<vsegment>
<ID>42</ID>
<points>32.5,-150.5,32.5,-148.5</points>
<connection>
<GID>98</GID>
<name>SEL_0</name></connection>
<intersection>-148.5 26</intersection></vsegment>
<vsegment>
<ID>43</ID>
<points>32.5,-137,32.5,-134.5</points>
<connection>
<GID>92</GID>
<name>SEL_0</name></connection>
<intersection>-134.5 19</intersection></vsegment>
<vsegment>
<ID>44</ID>
<points>33,-123,33,-121</points>
<connection>
<GID>86</GID>
<name>SEL_0</name></connection>
<intersection>-121 20</intersection></vsegment>
<vsegment>
<ID>45</ID>
<points>33,-109,33,-107</points>
<connection>
<GID>80</GID>
<name>SEL_0</name></connection>
<intersection>-107 21</intersection></vsegment>
<vsegment>
<ID>46</ID>
<points>33.5,-96,33.5,-93.5</points>
<connection>
<GID>74</GID>
<name>SEL_0</name></connection>
<intersection>-93.5 16</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>34,-81.5,34,-79</points>
<connection>
<GID>68</GID>
<name>SEL_0</name></connection>
<intersection>-79 11</intersection></vsegment>
<vsegment>
<ID>48</ID>
<points>34.5,-66.5,34.5,-64.5</points>
<connection>
<GID>62</GID>
<name>SEL_0</name></connection>
<intersection>-64.5 14</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>34.5,-50.5,34.5,-48.5</points>
<connection>
<GID>56</GID>
<name>SEL_0</name></connection>
<intersection>-48.5 15</intersection></vsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29.5,-22.5,33.5,-22.5</points>
<connection>
<GID>34</GID>
<name>IN_1</name></connection>
<connection>
<GID>37</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>32.5,-31.5,52.5,-31.5</points>
<intersection>32.5 5</intersection>
<intersection>52.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>52.5,-31.5,52.5,-23.5</points>
<intersection>-31.5 1</intersection>
<intersection>-23.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>49.5,-23.5,57,-23.5</points>
<connection>
<GID>35</GID>
<name>OUT_0</name></connection>
<connection>
<GID>39</GID>
<name>N_in0</name></connection>
<intersection>52.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>32.5,-31.5,32.5,-24.5</points>
<intersection>-31.5 1</intersection>
<intersection>-24.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>32.5,-24.5,33.5,-24.5</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<intersection>32.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>37,-38.5,43,-38.5</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<connection>
<GID>50</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29,-37.5,33,-37.5</points>
<connection>
<GID>52</GID>
<name>OUT_0</name></connection>
<connection>
<GID>50</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>32,-46.5,52,-46.5</points>
<intersection>32 5</intersection>
<intersection>52 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>52,-46.5,52,-38.5</points>
<intersection>-46.5 1</intersection>
<intersection>-38.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>49,-38.5,56.5,-38.5</points>
<connection>
<GID>53</GID>
<name>N_in0</name></connection>
<connection>
<GID>51</GID>
<name>OUT_0</name></connection>
<intersection>52 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>32,-46.5,32,-39.5</points>
<intersection>-46.5 1</intersection>
<intersection>-39.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>32,-39.5,33,-39.5</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>32 5</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>36.5,-53,42.5,-53</points>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<connection>
<GID>56</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-52,32.5,-52</points>
<connection>
<GID>56</GID>
<name>IN_1</name></connection>
<connection>
<GID>58</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-61,51.5,-61</points>
<intersection>31.5 5</intersection>
<intersection>51.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>51.5,-61,51.5,-53</points>
<intersection>-61 1</intersection>
<intersection>-53 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>48.5,-53,56,-53</points>
<connection>
<GID>59</GID>
<name>N_in0</name></connection>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection>
<intersection>51.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>31.5,-61,31.5,-54</points>
<intersection>-61 1</intersection>
<intersection>-54 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>31.5,-54,32.5,-54</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>31.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>36.5,-69,42.5,-69</points>
<connection>
<GID>62</GID>
<name>OUT</name></connection>
<connection>
<GID>63</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-68,32.5,-68</points>
<connection>
<GID>62</GID>
<name>IN_1</name></connection>
<connection>
<GID>64</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31.5,-77,51.5,-77</points>
<intersection>31.5 5</intersection>
<intersection>51.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>51.5,-77,51.5,-69</points>
<intersection>-77 1</intersection>
<intersection>-69 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>48.5,-69,56,-69</points>
<connection>
<GID>63</GID>
<name>OUT_0</name></connection>
<connection>
<GID>65</GID>
<name>N_in0</name></connection>
<intersection>51.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>31.5,-77,31.5,-70</points>
<intersection>-77 1</intersection>
<intersection>-70 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>31.5,-70,32.5,-70</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>31.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>36,-84,42,-84</points>
<connection>
<GID>68</GID>
<name>OUT</name></connection>
<connection>
<GID>69</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28,-83,32,-83</points>
<connection>
<GID>70</GID>
<name>OUT_0</name></connection>
<connection>
<GID>68</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31,-92,51,-92</points>
<intersection>31 5</intersection>
<intersection>51 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>51,-92,51,-84</points>
<intersection>-92 1</intersection>
<intersection>-84 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>48,-84,55.5,-84</points>
<connection>
<GID>69</GID>
<name>OUT_0</name></connection>
<connection>
<GID>71</GID>
<name>N_in0</name></connection>
<intersection>51 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>31,-92,31,-85</points>
<intersection>-92 1</intersection>
<intersection>-85 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>31,-85,32,-85</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<intersection>31 5</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35.5,-98.5,41.5,-98.5</points>
<connection>
<GID>75</GID>
<name>IN_0</name></connection>
<connection>
<GID>74</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27.5,-97.5,31.5,-97.5</points>
<connection>
<GID>76</GID>
<name>OUT_0</name></connection>
<connection>
<GID>74</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-106.5,50.5,-106.5</points>
<intersection>30.5 5</intersection>
<intersection>50.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>50.5,-106.5,50.5,-98.5</points>
<intersection>-106.5 1</intersection>
<intersection>-98.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>47.5,-98.5,55,-98.5</points>
<connection>
<GID>77</GID>
<name>N_in0</name></connection>
<connection>
<GID>75</GID>
<name>OUT_0</name></connection>
<intersection>50.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>30.5,-106.5,30.5,-99.5</points>
<intersection>-106.5 1</intersection>
<intersection>-99.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>30.5,-99.5,31.5,-99.5</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>30.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35,-111.5,41,-111.5</points>
<connection>
<GID>80</GID>
<name>OUT</name></connection>
<connection>
<GID>81</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27,-110.5,31,-110.5</points>
<connection>
<GID>82</GID>
<name>OUT_0</name></connection>
<connection>
<GID>80</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30,-119.5,50,-119.5</points>
<intersection>30 5</intersection>
<intersection>50 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>50,-119.5,50,-111.5</points>
<intersection>-119.5 1</intersection>
<intersection>-111.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>47,-111.5,54.5,-111.5</points>
<connection>
<GID>81</GID>
<name>OUT_0</name></connection>
<connection>
<GID>83</GID>
<name>N_in0</name></connection>
<intersection>50 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>30,-119.5,30,-112.5</points>
<intersection>-119.5 1</intersection>
<intersection>-112.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>30,-112.5,31,-112.5</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<intersection>30 5</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35,-125.5,41,-125.5</points>
<connection>
<GID>87</GID>
<name>IN_0</name></connection>
<connection>
<GID>86</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27,-124.5,31,-124.5</points>
<connection>
<GID>88</GID>
<name>OUT_0</name></connection>
<connection>
<GID>86</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30,-133.5,50,-133.5</points>
<intersection>30 5</intersection>
<intersection>50 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>50,-133.5,50,-125.5</points>
<intersection>-133.5 1</intersection>
<intersection>-125.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>47,-125.5,54.5,-125.5</points>
<connection>
<GID>89</GID>
<name>N_in0</name></connection>
<connection>
<GID>87</GID>
<name>OUT_0</name></connection>
<intersection>50 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>30,-133.5,30,-126.5</points>
<intersection>-133.5 1</intersection>
<intersection>-126.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>30,-126.5,31,-126.5</points>
<connection>
<GID>86</GID>
<name>IN_0</name></connection>
<intersection>30 5</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34.5,-139.5,40.5,-139.5</points>
<connection>
<GID>93</GID>
<name>IN_0</name></connection>
<connection>
<GID>92</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-138.5,30.5,-138.5</points>
<connection>
<GID>94</GID>
<name>OUT_0</name></connection>
<connection>
<GID>92</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29.5,-147.5,49.5,-147.5</points>
<intersection>29.5 5</intersection>
<intersection>49.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>49.5,-147.5,49.5,-139.5</points>
<intersection>-147.5 1</intersection>
<intersection>-139.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>46.5,-139.5,54,-139.5</points>
<connection>
<GID>95</GID>
<name>N_in0</name></connection>
<connection>
<GID>93</GID>
<name>OUT_0</name></connection>
<intersection>49.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>29.5,-147.5,29.5,-140.5</points>
<intersection>-147.5 1</intersection>
<intersection>-140.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>29.5,-140.5,30.5,-140.5</points>
<connection>
<GID>92</GID>
<name>IN_0</name></connection>
<intersection>29.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34.5,-153,40.5,-153</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<connection>
<GID>98</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-152,30.5,-152</points>
<connection>
<GID>100</GID>
<name>OUT_0</name></connection>
<connection>
<GID>98</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29.5,-161,49.5,-161</points>
<intersection>29.5 5</intersection>
<intersection>49.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>49.5,-161,49.5,-153</points>
<intersection>-161 1</intersection>
<intersection>-153 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>46.5,-153,54,-153</points>
<connection>
<GID>101</GID>
<name>N_in0</name></connection>
<connection>
<GID>99</GID>
<name>OUT_0</name></connection>
<intersection>49.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>29.5,-161,29.5,-154</points>
<intersection>-161 1</intersection>
<intersection>-154 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>29.5,-154,30.5,-154</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>29.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35,-169,41,-169</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<connection>
<GID>104</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27,-168,31,-168</points>
<connection>
<GID>106</GID>
<name>OUT_0</name></connection>
<connection>
<GID>104</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30,-177,50,-177</points>
<intersection>30 5</intersection>
<intersection>50 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>50,-177,50,-169</points>
<intersection>-177 1</intersection>
<intersection>-169 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>47,-169,54.5,-169</points>
<connection>
<GID>107</GID>
<name>N_in0</name></connection>
<connection>
<GID>105</GID>
<name>OUT_0</name></connection>
<intersection>50 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>30,-177,30,-170</points>
<intersection>-177 1</intersection>
<intersection>-170 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>30,-170,31,-170</points>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<intersection>30 5</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34.5,-183.5,40.5,-183.5</points>
<connection>
<GID>110</GID>
<name>OUT</name></connection>
<connection>
<GID>111</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-182.5,30.5,-182.5</points>
<connection>
<GID>112</GID>
<name>OUT_0</name></connection>
<connection>
<GID>110</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29.5,-191.5,49.5,-191.5</points>
<intersection>29.5 5</intersection>
<intersection>49.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>49.5,-191.5,49.5,-183.5</points>
<intersection>-191.5 1</intersection>
<intersection>-183.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>46.5,-183.5,54,-183.5</points>
<connection>
<GID>113</GID>
<name>N_in0</name></connection>
<connection>
<GID>111</GID>
<name>OUT_0</name></connection>
<intersection>49.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>29.5,-191.5,29.5,-184.5</points>
<intersection>-191.5 1</intersection>
<intersection>-184.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>29.5,-184.5,30.5,-184.5</points>
<connection>
<GID>110</GID>
<name>IN_0</name></connection>
<intersection>29.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>54</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34.5,-199.5,40.5,-199.5</points>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<connection>
<GID>116</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-198.5,30.5,-198.5</points>
<connection>
<GID>118</GID>
<name>OUT_0</name></connection>
<connection>
<GID>116</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29.5,-207.5,49.5,-207.5</points>
<intersection>29.5 5</intersection>
<intersection>49.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>49.5,-207.5,49.5,-199.5</points>
<intersection>-207.5 1</intersection>
<intersection>-199.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>46.5,-199.5,54,-199.5</points>
<connection>
<GID>119</GID>
<name>N_in0</name></connection>
<connection>
<GID>117</GID>
<name>OUT_0</name></connection>
<intersection>49.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>29.5,-207.5,29.5,-200.5</points>
<intersection>-207.5 1</intersection>
<intersection>-200.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>29.5,-200.5,30.5,-200.5</points>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<intersection>29.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>32.5,-215.5,38.5,-215.5</points>
<connection>
<GID>122</GID>
<name>OUT</name></connection>
<connection>
<GID>123</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>24.5,-214.5,28.5,-214.5</points>
<connection>
<GID>124</GID>
<name>OUT_0</name></connection>
<connection>
<GID>122</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27.5,-223.5,47.5,-223.5</points>
<intersection>27.5 5</intersection>
<intersection>47.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>47.5,-223.5,47.5,-215.5</points>
<intersection>-223.5 1</intersection>
<intersection>-215.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>44.5,-215.5,52,-215.5</points>
<connection>
<GID>123</GID>
<name>OUT_0</name></connection>
<connection>
<GID>125</GID>
<name>N_in0</name></connection>
<intersection>47.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>27.5,-223.5,27.5,-216.5</points>
<intersection>-223.5 1</intersection>
<intersection>-216.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>27.5,-216.5,28.5,-216.5</points>
<connection>
<GID>122</GID>
<name>IN_0</name></connection>
<intersection>27.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-232,40,-232</points>
<connection>
<GID>129</GID>
<name>IN_0</name></connection>
<connection>
<GID>128</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26,-231,30,-231</points>
<connection>
<GID>130</GID>
<name>OUT_0</name></connection>
<connection>
<GID>128</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29,-240,49,-240</points>
<intersection>29 5</intersection>
<intersection>49 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>49,-240,49,-232</points>
<intersection>-240 1</intersection>
<intersection>-232 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>46,-232,53.5,-232</points>
<connection>
<GID>131</GID>
<name>N_in0</name></connection>
<connection>
<GID>129</GID>
<name>OUT_0</name></connection>
<intersection>49 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>29,-240,29,-233</points>
<intersection>-240 1</intersection>
<intersection>-233 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>29,-233,30,-233</points>
<connection>
<GID>128</GID>
<name>IN_0</name></connection>
<intersection>29 5</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33,-248,39,-248</points>
<connection>
<GID>135</GID>
<name>IN_0</name></connection>
<connection>
<GID>134</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25,-247,29,-247</points>
<connection>
<GID>136</GID>
<name>OUT_0</name></connection>
<connection>
<GID>134</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28,-256,48,-256</points>
<intersection>28 5</intersection>
<intersection>48 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>48,-256,48,-248</points>
<intersection>-256 1</intersection>
<intersection>-248 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>45,-248,52.5,-248</points>
<connection>
<GID>137</GID>
<name>N_in0</name></connection>
<connection>
<GID>135</GID>
<name>OUT_0</name></connection>
<intersection>48 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>28,-256,28,-249</points>
<intersection>-256 1</intersection>
<intersection>-249 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>28,-249,29,-249</points>
<connection>
<GID>134</GID>
<name>IN_0</name></connection>
<intersection>28 5</intersection></hsegment></shape></wire>
<wire>
<ID>66</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-263,40,-263</points>
<connection>
<GID>140</GID>
<name>OUT</name></connection>
<connection>
<GID>141</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>67</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26,-262,30,-262</points>
<connection>
<GID>142</GID>
<name>OUT_0</name></connection>
<connection>
<GID>140</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>29,-271,49,-271</points>
<intersection>29 5</intersection>
<intersection>49 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>49,-271,49,-263</points>
<intersection>-271 1</intersection>
<intersection>-263 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>46,-263,53.5,-263</points>
<connection>
<GID>141</GID>
<name>OUT_0</name></connection>
<connection>
<GID>143</GID>
<name>N_in0</name></connection>
<intersection>49 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>29,-271,29,-264</points>
<intersection>-271 1</intersection>
<intersection>-264 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>29,-264,30,-264</points>
<connection>
<GID>140</GID>
<name>IN_0</name></connection>
<intersection>29 5</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8.5,-266,8.5,-26.5</points>
<intersection>-266 24</intersection>
<intersection>-251 25</intersection>
<intersection>-235 22</intersection>
<intersection>-218.5 19</intersection>
<intersection>-202.5 21</intersection>
<intersection>-186.5 15</intersection>
<intersection>-172 16</intersection>
<intersection>-156 13</intersection>
<intersection>-147 1</intersection>
<intersection>-128.5 17</intersection>
<intersection>-114.5 8</intersection>
<intersection>-101.5 10</intersection>
<intersection>-87 6</intersection>
<intersection>-72 9</intersection>
<intersection>-56 4</intersection>
<intersection>-41.5 11</intersection>
<intersection>-26.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>1,-147,8.5,-147</points>
<connection>
<GID>38</GID>
<name>CLK</name></connection>
<intersection>8.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>8.5,-26.5,43.5,-26.5</points>
<connection>
<GID>35</GID>
<name>clock</name></connection>
<intersection>8.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>8.5,-56,42.5,-56</points>
<connection>
<GID>57</GID>
<name>clock</name></connection>
<intersection>8.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>8.5,-87,42,-87</points>
<connection>
<GID>69</GID>
<name>clock</name></connection>
<intersection>8.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>8.5,-114.5,41,-114.5</points>
<connection>
<GID>81</GID>
<name>clock</name></connection>
<intersection>8.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>8.5,-72,42.5,-72</points>
<connection>
<GID>63</GID>
<name>clock</name></connection>
<intersection>8.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>8.5,-101.5,41.5,-101.5</points>
<connection>
<GID>75</GID>
<name>clock</name></connection>
<intersection>8.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>8.5,-41.5,43,-41.5</points>
<connection>
<GID>51</GID>
<name>clock</name></connection>
<intersection>8.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>8.5,-156,40.5,-156</points>
<connection>
<GID>99</GID>
<name>clock</name></connection>
<intersection>8.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>8.5,-186.5,40.5,-186.5</points>
<connection>
<GID>111</GID>
<name>clock</name></connection>
<intersection>8.5 0</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>8.5,-172,41,-172</points>
<connection>
<GID>105</GID>
<name>clock</name></connection>
<intersection>8.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>8.5,-128.5,41,-128.5</points>
<connection>
<GID>87</GID>
<name>clock</name></connection>
<intersection>8.5 0</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>8.5,-218.5,38.5,-218.5</points>
<connection>
<GID>123</GID>
<name>clock</name></connection>
<intersection>8.5 0</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>8.5,-202.5,40.5,-202.5</points>
<connection>
<GID>117</GID>
<name>clock</name></connection>
<intersection>8.5 0</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>8.5,-235,40,-235</points>
<connection>
<GID>129</GID>
<name>clock</name></connection>
<intersection>8.5 0</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>8.5,-266,40,-266</points>
<connection>
<GID>141</GID>
<name>clock</name></connection>
<intersection>8.5 0</intersection></hsegment>
<hsegment>
<ID>25</ID>
<points>8.5,-251,39,-251</points>
<connection>
<GID>135</GID>
<name>clock</name></connection>
<intersection>8.5 0</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>-50.8003,59.2835,134.675,-34.1197</PageViewport>
<gate>
<ID>146</ID>
<type>AA_TOGGLE</type>
<position>29,23</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>147</ID>
<type>AA_TOGGLE</type>
<position>29,20</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>148</ID>
<type>AA_TOGGLE</type>
<position>29,17</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>149</ID>
<type>AA_TOGGLE</type>
<position>29,14</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>150</ID>
<type>AA_TOGGLE</type>
<position>29,11</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>151</ID>
<type>AA_TOGGLE</type>
<position>29,8</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>152</ID>
<type>AA_TOGGLE</type>
<position>29,5</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>153</ID>
<type>AA_TOGGLE</type>
<position>29,2</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>154</ID>
<type>AA_TOGGLE</type>
<position>29,-1</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>155</ID>
<type>AA_TOGGLE</type>
<position>29,-4</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>156</ID>
<type>AA_TOGGLE</type>
<position>29,-7</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>157</ID>
<type>AA_TOGGLE</type>
<position>29,-10</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>158</ID>
<type>AA_TOGGLE</type>
<position>29,-13</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>159</ID>
<type>AA_TOGGLE</type>
<position>29,-16</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>160</ID>
<type>AA_TOGGLE</type>
<position>29,-19</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>161</ID>
<type>AA_TOGGLE</type>
<position>29,-22</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate></page 2>
<page 3>
<PageViewport>0,37.7538,439.646,-183.646</PageViewport></page 3>
<page 4>
<PageViewport>0,37.7538,439.646,-183.646</PageViewport></page 4>
<page 5>
<PageViewport>0,37.7538,439.646,-183.646</PageViewport></page 5>
<page 6>
<PageViewport>0,37.7538,439.646,-183.646</PageViewport></page 6>
<page 7>
<PageViewport>0,37.7538,439.646,-183.646</PageViewport></page 7>
<page 8>
<PageViewport>0,37.7538,439.646,-183.646</PageViewport></page 8>
<page 9>
<PageViewport>0,37.7538,439.646,-183.646</PageViewport></page 9></circuit>