<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-11.4,8.66667,174.467,-84.9333</PageViewport>
<gate>
<ID>11</ID>
<type>AA_TOGGLE</type>
<position>19,-4</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>13</ID>
<type>AA_TOGGLE</type>
<position>32.5,-4</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_TOGGLE</type>
<position>45.5,-4</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_TOGGLE</type>
<position>51.5,-4</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>19</ID>
<type>AA_TOGGLE</type>
<position>57.5,-4</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_TOGGLE</type>
<position>63.5,-4</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_TOGGLE</type>
<position>6,-23</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_TOGGLE</type>
<position>6,-31</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_LABEL</type>
<position>19.5,0</position>
<gparam>LABEL_TEXT zx</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>AA_LABEL</type>
<position>33,0</position>
<gparam>LABEL_TEXT nx</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>AA_LABEL</type>
<position>45.5,0</position>
<gparam>LABEL_TEXT zy</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>31</ID>
<type>AA_LABEL</type>
<position>51.5,0</position>
<gparam>LABEL_TEXT ny</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>33</ID>
<type>AA_LABEL</type>
<position>57.5,-0.5</position>
<gparam>LABEL_TEXT f</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>AA_LABEL</type>
<position>63.5,-0.5</position>
<gparam>LABEL_TEXT no</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>37</ID>
<type>AA_LABEL</type>
<position>3,-22</position>
<gparam>LABEL_TEXT x</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>AA_LABEL</type>
<position>3,-30.5</position>
<gparam>LABEL_TEXT y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>43</ID>
<type>AA_INVERTER</type>
<position>25.5,-4</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>45</ID>
<type>AA_AND2</type>
<position>33,-19</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>47</ID>
<type>GA_LED</type>
<position>40.5,-19</position>
<input>
<ID>N_in0</ID>4 </input>
<input>
<ID>N_in1</ID>4 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>49</ID>
<type>AA_LABEL</type>
<position>19.5,-12.5</position>
<gparam>LABEL_TEXT if zx then make x be zero</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>56</ID>
<type>AA_LABEL</type>
<position>51,-22.5</position>
<gparam>LABEL_TEXT if nx then negate x</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>58</ID>
<type>AA_INVERTER</type>
<position>25,-29</position>
<input>
<ID>IN_0</ID>3 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>60</ID>
<type>AA_INVERTER</type>
<position>25,-34</position>
<input>
<ID>IN_0</ID>3 </input>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>62</ID>
<type>AA_INVERTER</type>
<position>39,-4</position>
<input>
<ID>IN_0</ID>8 </input>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>64</ID>
<type>AA_AND2</type>
<position>46.5,-28</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>66</ID>
<type>AA_AND2</type>
<position>46.5,-33</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>13 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>68</ID>
<type>AE_OR2</type>
<position>55.5,-30.5</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>15 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>70</ID>
<type>GA_LED</type>
<position>61.5,-30.5</position>
<input>
<ID>N_in0</ID>16 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21,-4,22.5,-4</points>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection>
<connection>
<GID>43</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-4,30,-4</points>
<connection>
<GID>43</GID>
<name>OUT_0</name></connection>
<intersection>30 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>30,-18,30,-4</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>-4 1</intersection></vsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19.5,-34,19.5,-20</points>
<intersection>-34 5</intersection>
<intersection>-29 3</intersection>
<intersection>-23 1</intersection>
<intersection>-20 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8,-23,19.5,-23</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<intersection>19.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>19.5,-20,30,-20</points>
<connection>
<GID>45</GID>
<name>IN_1</name></connection>
<intersection>19.5 0</intersection>
<intersection>30 6</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>19.5,-29,22,-29</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>19.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>19.5,-34,22,-34</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>19.5 0</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>30,-29,30,-20</points>
<intersection>-29 7</intersection>
<intersection>-20 2</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>30,-29,43.5,-29</points>
<connection>
<GID>64</GID>
<name>IN_1</name></connection>
<intersection>30 6</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>36,-19,41.5,-19</points>
<connection>
<GID>47</GID>
<name>N_in1</name></connection>
<connection>
<GID>45</GID>
<name>OUT</name></connection>
<connection>
<GID>47</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34.5,-4,36,-4</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<connection>
<GID>13</GID>
<name>OUT_0</name></connection>
<intersection>36 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>36,-32,36,-4</points>
<intersection>-32 4</intersection>
<intersection>-4 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>36,-32,43.5,-32</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>36 3</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,-27,42.5,-4</points>
<intersection>-27 4</intersection>
<intersection>-4 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>42,-4,42.5,-4</points>
<connection>
<GID>62</GID>
<name>OUT_0</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>42.5,-27,43.5,-27</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<intersection>42.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28,-34,43.5,-34</points>
<connection>
<GID>60</GID>
<name>OUT_0</name></connection>
<connection>
<GID>66</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-29.5,51,-28</points>
<intersection>-29.5 1</intersection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51,-29.5,52.5,-29.5</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<intersection>51 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49.5,-28,51,-28</points>
<connection>
<GID>64</GID>
<name>OUT</name></connection>
<intersection>51 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-33,51,-31.5</points>
<intersection>-33 2</intersection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51,-31.5,52.5,-31.5</points>
<connection>
<GID>68</GID>
<name>IN_1</name></connection>
<intersection>51 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49.5,-33,51,-33</points>
<connection>
<GID>66</GID>
<name>OUT</name></connection>
<intersection>51 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58.5,-30.5,60.5,-30.5</points>
<connection>
<GID>70</GID>
<name>N_in0</name></connection>
<connection>
<GID>68</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 1>
<page 2>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 2>
<page 3>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 3>
<page 4>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 4>
<page 5>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 5>
<page 6>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 6>
<page 7>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 7>
<page 8>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 8>
<page 9>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 9></circuit>