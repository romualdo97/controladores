<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>30.4937,-15.3562,108.906,-54.8438</PageViewport>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>42.5,-21</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>37,-21</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>6</ID>
<type>AI_XOR2</type>
<position>51,-28</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_LABEL</type>
<position>42.5,-17.5</position>
<gparam>LABEL_TEXT a</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>9</ID>
<type>AA_LABEL</type>
<position>37,-17.5</position>
<gparam>LABEL_TEXT b</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>11</ID>
<type>AA_LABEL</type>
<position>64,-27.5</position>
<gparam>LABEL_TEXT sum</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>13</ID>
<type>AA_AND2</type>
<position>51,-36.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>15</ID>
<type>AA_LABEL</type>
<position>64.5,-35.5</position>
<gparam>LABEL_TEXT carry</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>17</ID>
<type>GA_LED</type>
<position>56.5,-28</position>
<input>
<ID>N_in0</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>GA_LED</type>
<position>56.5,-36.5</position>
<input>
<ID>N_in0</ID>4 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-35.5,45,-21</points>
<intersection>-35.5 9</intersection>
<intersection>-27 2</intersection>
<intersection>-21 7</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>45,-27,48,-27</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>44.5,-21,45,-21</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>45,-35.5,48,-35.5</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-37.5,40,-21</points>
<intersection>-37.5 4</intersection>
<intersection>-29 2</intersection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39,-21,40,-21</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>40 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>40,-29,48,-29</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>40 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>40,-37.5,48,-37.5</points>
<connection>
<GID>13</GID>
<name>IN_1</name></connection>
<intersection>40 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54,-28,55.5,-28</points>
<connection>
<GID>17</GID>
<name>N_in0</name></connection>
<connection>
<GID>6</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54,-36.5,55.5,-36.5</points>
<connection>
<GID>19</GID>
<name>N_in0</name></connection>
<connection>
<GID>13</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 1>
<page 2>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 2>
<page 3>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 3>
<page 4>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 4>
<page 5>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 5>
<page 6>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 6>
<page 7>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 7>
<page 8>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 8>
<page 9>
<PageViewport>0,0,139.4,-70.2</PageViewport></page 9></circuit>