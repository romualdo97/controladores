<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-31.063,76.6229,652.896,-267.81</PageViewport>
<gate>
<ID>2</ID>
<type>AA_INVERTER</type>
<position>25.5,-42.5</position>
<input>
<ID>IN_0</ID>5 </input>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_INVERTER</type>
<position>40.5,-42.5</position>
<input>
<ID>IN_0</ID>6 </input>
<output>
<ID>OUT_0</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>5</ID>
<type>AA_AND2</type>
<position>31.5,-57</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>30 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>GA_LED</type>
<position>39,-57</position>
<input>
<ID>N_in0</ID>9 </input>
<input>
<ID>N_in1</ID>9 </input>
<input>
<ID>N_in2</ID>9 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>7</ID>
<type>AA_LABEL</type>
<position>18,-50.5</position>
<gparam>LABEL_TEXT if zy then make y be zero</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>AA_LABEL</type>
<position>49.5,-60.5</position>
<gparam>LABEL_TEXT if ny then negate y</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>9</ID>
<type>AA_INVERTER</type>
<position>25.5,-72</position>
<input>
<ID>IN_0</ID>30 </input>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_AND2</type>
<position>46.5,-66</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>30 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>11</ID>
<type>AA_TOGGLE</type>
<position>19,-4</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_AND2</type>
<position>45,-71</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>13</ID>
<type>AA_TOGGLE</type>
<position>32.5,-4</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>14</ID>
<type>AE_OR2</type>
<position>54,-68.5</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>17 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>15</ID>
<type>GA_LED</type>
<position>60,-68.5</position>
<input>
<ID>N_in0</ID>18 </input>
<input>
<ID>N_in1</ID>37 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>17</ID>
<type>AA_TOGGLE</type>
<position>18.5,-42.5</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_TOGGLE</type>
<position>33,-42.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>19</ID>
<type>AA_TOGGLE</type>
<position>92,-2.5</position>
<output>
<ID>OUT_0</ID>52 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_TOGGLE</type>
<position>105.5,-2.5</position>
<output>
<ID>OUT_0</ID>57 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_TOGGLE</type>
<position>6,-23</position>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>23</ID>
<type>AA_LABEL</type>
<position>100.5,-50</position>
<gparam>LABEL_TEXT if f then x+y else x&y</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>AA_TOGGLE</type>
<position>6,-58</position>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_LABEL</type>
<position>19.5,0</position>
<gparam>LABEL_TEXT zx</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>AA_LABEL</type>
<position>33,0</position>
<gparam>LABEL_TEXT nx</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>AA_LABEL</type>
<position>19,-38.5</position>
<gparam>LABEL_TEXT zy</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>31</ID>
<type>AA_LABEL</type>
<position>33.5,-38.5</position>
<gparam>LABEL_TEXT ny</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>33</ID>
<type>AA_LABEL</type>
<position>92,1.5</position>
<gparam>LABEL_TEXT f</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>AA_LABEL</type>
<position>105.5,1</position>
<gparam>LABEL_TEXT no</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>37</ID>
<type>AA_LABEL</type>
<position>3,-22</position>
<gparam>LABEL_TEXT x</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>AA_LABEL</type>
<position>3,-57.5</position>
<gparam>LABEL_TEXT y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>GA_LED</type>
<position>88.5,-54</position>
<input>
<ID>N_in0</ID>43 </input>
<input>
<ID>N_in1</ID>51 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>43</ID>
<type>AA_INVERTER</type>
<position>25.5,-4</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>45</ID>
<type>AA_AND2</type>
<position>33,-19</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>28 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>47</ID>
<type>GA_LED</type>
<position>40.5,-19</position>
<input>
<ID>N_in0</ID>4 </input>
<input>
<ID>N_in1</ID>4 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>49</ID>
<type>AA_LABEL</type>
<position>19.5,-12.5</position>
<gparam>LABEL_TEXT if zx then make x be zero</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>54</ID>
<type>AA_FULLADDER_1BIT</type>
<position>81,-54</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_B_0</ID>37 </input>
<output>
<ID>OUT_0</ID>43 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>56</ID>
<type>AA_LABEL</type>
<position>51,-22.5</position>
<gparam>LABEL_TEXT if nx then negate x</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>AA_INVERTER</type>
<position>25,-34</position>
<input>
<ID>IN_0</ID>28 </input>
<output>
<ID>OUT_0</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>62</ID>
<type>AA_INVERTER</type>
<position>39,-4</position>
<input>
<ID>IN_0</ID>8 </input>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>64</ID>
<type>AA_AND2</type>
<position>46.5,-28</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>28 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>66</ID>
<type>AA_AND2</type>
<position>46.5,-33</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>31 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>67</ID>
<type>GA_LED</type>
<position>135.5,-45.5</position>
<input>
<ID>N_in0</ID>56 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>68</ID>
<type>AE_OR2</type>
<position>55.5,-30.5</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>15 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>70</ID>
<type>GA_LED</type>
<position>61.5,-30.5</position>
<input>
<ID>N_in0</ID>16 </input>
<input>
<ID>N_in1</ID>36 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>73</ID>
<type>AA_AND2</type>
<position>79.5,-38</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>37 </input>
<output>
<ID>OUT</ID>47 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>75</ID>
<type>GA_LED</type>
<position>86,-38</position>
<input>
<ID>N_in0</ID>47 </input>
<input>
<ID>N_in1</ID>50 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>76</ID>
<type>AA_LABEL</type>
<position>83,-48.5</position>
<gparam>LABEL_TEXT xo plus yo</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>77</ID>
<type>AA_LABEL</type>
<position>82,-33</position>
<gparam>LABEL_TEXT xo and yo</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>79</ID>
<type>AA_MUX_2x1</type>
<position>97.5,-46</position>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>50 </input>
<output>
<ID>OUT</ID>58 </output>
<input>
<ID>SEL_0</ID>52 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>81</ID>
<type>AA_MUX_2x1</type>
<position>120.5,-45.5</position>
<input>
<ID>IN_0</ID>59 </input>
<input>
<ID>IN_1</ID>55 </input>
<output>
<ID>OUT</ID>56 </output>
<input>
<ID>SEL_0</ID>57 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>83</ID>
<type>AA_INVERTER</type>
<position>108.5,-41</position>
<input>
<ID>IN_0</ID>59 </input>
<output>
<ID>OUT_0</ID>55 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>85</ID>
<type>GA_LED</type>
<position>102.5,-46</position>
<input>
<ID>N_in0</ID>58 </input>
<input>
<ID>N_in1</ID>59 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>21,-4,22.5,-4</points>
<connection>
<GID>11</GID>
<name>OUT_0</name></connection>
<connection>
<GID>43</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-4,30,-4</points>
<connection>
<GID>43</GID>
<name>OUT_0</name></connection>
<intersection>30 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>30,-18,30,-4</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>-4 1</intersection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>36,-19,41.5,-19</points>
<connection>
<GID>47</GID>
<name>N_in1</name></connection>
<connection>
<GID>45</GID>
<name>OUT</name></connection>
<connection>
<GID>47</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20.5,-42.5,22.5,-42.5</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<connection>
<GID>17</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35,-42.5,37.5,-42.5</points>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>35.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>35.5,-70,35.5,-42.5</points>
<intersection>-70 4</intersection>
<intersection>-42.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>35.5,-70,42,-70</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>35.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34.5,-4,36,-4</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<connection>
<GID>13</GID>
<name>OUT_0</name></connection>
<intersection>36 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>36,-32,36,-4</points>
<intersection>-32 4</intersection>
<intersection>-4 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>36,-32,43.5,-32</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>36 3</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34.5,-57,40,-57</points>
<connection>
<GID>6</GID>
<name>N_in1</name></connection>
<connection>
<GID>6</GID>
<name>N_in0</name></connection>
<connection>
<GID>5</GID>
<name>OUT</name></connection>
<intersection>39 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>39,-58,39,-57</points>
<connection>
<GID>6</GID>
<name>N_in2</name></connection>
<intersection>-57 1</intersection></vsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28.5,-72,42,-72</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<connection>
<GID>9</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-67.5,49.5,-66</points>
<connection>
<GID>10</GID>
<name>OUT</name></connection>
<intersection>-67.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49.5,-67.5,51,-67.5</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,-27,42.5,-4</points>
<intersection>-27 4</intersection>
<intersection>-4 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>42,-4,42.5,-4</points>
<connection>
<GID>62</GID>
<name>OUT_0</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>42.5,-27,43.5,-27</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<intersection>42.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-29.5,51,-28</points>
<intersection>-29.5 1</intersection>
<intersection>-28 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51,-29.5,52.5,-29.5</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<intersection>51 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49.5,-28,51,-28</points>
<connection>
<GID>64</GID>
<name>OUT</name></connection>
<intersection>51 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-33,51,-31.5</points>
<intersection>-33 2</intersection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>51,-31.5,52.5,-31.5</points>
<connection>
<GID>68</GID>
<name>IN_1</name></connection>
<intersection>51 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>49.5,-33,51,-33</points>
<connection>
<GID>66</GID>
<name>OUT</name></connection>
<intersection>51 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58.5,-30.5,60.5,-30.5</points>
<connection>
<GID>70</GID>
<name>N_in0</name></connection>
<connection>
<GID>68</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>49.5,-71,49.5,-69.5</points>
<intersection>-71 2</intersection>
<intersection>-69.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>49.5,-69.5,51,-69.5</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>49.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>48,-71,49.5,-71</points>
<connection>
<GID>12</GID>
<name>OUT</name></connection>
<intersection>49.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-68.5,59,-68.5</points>
<connection>
<GID>14</GID>
<name>OUT</name></connection>
<connection>
<GID>15</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-56,28.5,-42.5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<connection>
<GID>5</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-65,43.5,-42.5</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<connection>
<GID>10</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>19,-34,19,-20</points>
<intersection>-34 5</intersection>
<intersection>-29 4</intersection>
<intersection>-23 1</intersection>
<intersection>-20 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8,-23,19,-23</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<intersection>19 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>19,-20,30,-20</points>
<connection>
<GID>45</GID>
<name>IN_1</name></connection>
<intersection>19 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>19,-29,43.5,-29</points>
<connection>
<GID>64</GID>
<name>IN_1</name></connection>
<intersection>19 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>19,-34,22,-34</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>19 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>8,-58,28.5,-58</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<connection>
<GID>5</GID>
<name>IN_1</name></connection>
<intersection>20.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>20.5,-72,20.5,-58</points>
<intersection>-72 6</intersection>
<intersection>-67 5</intersection>
<intersection>-58 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>20.5,-67,43.5,-67</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<intersection>20.5 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>20.5,-72,22.5,-72</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<intersection>20.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>28,-34,43.5,-34</points>
<connection>
<GID>60</GID>
<name>OUT_0</name></connection>
<connection>
<GID>66</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68,-53,68,-30.5</points>
<intersection>-53 1</intersection>
<intersection>-37 4</intersection>
<intersection>-30.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68,-53,78,-53</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>68 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>62.5,-30.5,68,-30.5</points>
<connection>
<GID>70</GID>
<name>N_in1</name></connection>
<intersection>68 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>68,-37,76.5,-37</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>68 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68,-68.5,68,-55</points>
<intersection>-68.5 2</intersection>
<intersection>-65.5 3</intersection>
<intersection>-55 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68,-55,78,-55</points>
<connection>
<GID>54</GID>
<name>IN_B_0</name></connection>
<intersection>68 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>61,-68.5,68,-68.5</points>
<connection>
<GID>15</GID>
<name>N_in1</name></connection>
<intersection>68 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>68,-65.5,76,-65.5</points>
<intersection>68 0</intersection>
<intersection>76 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>76,-65.5,76,-39</points>
<intersection>-65.5 3</intersection>
<intersection>-39 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>76,-39,76.5,-39</points>
<connection>
<GID>73</GID>
<name>IN_1</name></connection>
<intersection>76 6</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>84,-54,87.5,-54</points>
<connection>
<GID>42</GID>
<name>N_in0</name></connection>
<connection>
<GID>54</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82.5,-38,85,-38</points>
<connection>
<GID>73</GID>
<name>OUT</name></connection>
<connection>
<GID>75</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>91,-45,91,-38</points>
<intersection>-45 2</intersection>
<intersection>-38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>87,-38,91,-38</points>
<connection>
<GID>75</GID>
<name>N_in1</name></connection>
<intersection>91 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>91,-45,95.5,-45</points>
<connection>
<GID>79</GID>
<name>IN_1</name></connection>
<intersection>91 0</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92.5,-54,92.5,-47</points>
<intersection>-54 1</intersection>
<intersection>-47 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>89.5,-54,92.5,-54</points>
<connection>
<GID>42</GID>
<name>N_in1</name></connection>
<intersection>92.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>92.5,-47,95.5,-47</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>92.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97.5,-43.5,97.5,-2.5</points>
<connection>
<GID>79</GID>
<name>SEL_0</name></connection>
<intersection>-2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>94,-2.5,97.5,-2.5</points>
<connection>
<GID>19</GID>
<name>OUT_0</name></connection>
<intersection>97.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112.5,-44.5,112.5,-41</points>
<intersection>-44.5 1</intersection>
<intersection>-41 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>112.5,-44.5,118.5,-44.5</points>
<connection>
<GID>81</GID>
<name>IN_1</name></connection>
<intersection>112.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>111.5,-41,112.5,-41</points>
<connection>
<GID>83</GID>
<name>OUT_0</name></connection>
<intersection>112.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>122.5,-45.5,134.5,-45.5</points>
<connection>
<GID>67</GID>
<name>N_in0</name></connection>
<connection>
<GID>81</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>120.5,-43,120.5,-2.5</points>
<connection>
<GID>81</GID>
<name>SEL_0</name></connection>
<intersection>-2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107.5,-2.5,120.5,-2.5</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>120.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>99.5,-46,101.5,-46</points>
<connection>
<GID>85</GID>
<name>N_in0</name></connection>
<connection>
<GID>79</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-46.5,104.5,-41</points>
<intersection>-46.5 3</intersection>
<intersection>-46 1</intersection>
<intersection>-41 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>103.5,-46,104.5,-46</points>
<connection>
<GID>85</GID>
<name>N_in1</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104.5,-41,105.5,-41</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>104.5,-46.5,118.5,-46.5</points>
<connection>
<GID>81</GID>
<name>IN_0</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>116.039,-2.76362,532.482,-212.479</PageViewport>
<gate>
<ID>90</ID>
<type>AA_LABEL</type>
<position>69,-88</position>
<gparam>LABEL_TEXT if zy then make y be zero</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>91</ID>
<type>AA_LABEL</type>
<position>96.5,-87.5</position>
<gparam>LABEL_TEXT if ny then negate zyo</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>94</ID>
<type>AA_TOGGLE</type>
<position>69.5,-30</position>
<output>
<ID>OUT_0</ID>99 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>96</ID>
<type>AA_TOGGLE</type>
<position>88.5,-30</position>
<output>
<ID>OUT_0</ID>130 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>99</ID>
<type>AA_TOGGLE</type>
<position>69,-68.5</position>
<output>
<ID>OUT_0</ID>108 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>100</ID>
<type>AA_TOGGLE</type>
<position>83.5,-68.5</position>
<output>
<ID>OUT_0</ID>134 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>101</ID>
<type>AA_TOGGLE</type>
<position>142.5,-28.5</position>
<output>
<ID>OUT_0</ID>86 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>102</ID>
<type>AA_TOGGLE</type>
<position>156,-28.5</position>
<output>
<ID>OUT_0</ID>89 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>103</ID>
<type>AA_TOGGLE</type>
<position>56.5,-51</position>
<output>
<ID>OUT_0</ID>100 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>104</ID>
<type>AA_LABEL</type>
<position>152.5,-76</position>
<gparam>LABEL_TEXT if f then xo+yo else xo&yo</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>105</ID>
<type>AA_TOGGLE</type>
<position>56.5,-84</position>
<output>
<ID>OUT_0</ID>105 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>106</ID>
<type>AA_LABEL</type>
<position>70,-26</position>
<gparam>LABEL_TEXT zx</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>107</ID>
<type>AA_LABEL</type>
<position>89,-26</position>
<gparam>LABEL_TEXT nx</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>108</ID>
<type>AA_LABEL</type>
<position>69.5,-64.5</position>
<gparam>LABEL_TEXT zy</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>109</ID>
<type>AA_LABEL</type>
<position>84,-64.5</position>
<gparam>LABEL_TEXT ny</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>110</ID>
<type>AA_LABEL</type>
<position>142.5,-24.5</position>
<gparam>LABEL_TEXT f</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>111</ID>
<type>AA_LABEL</type>
<position>156,-25</position>
<gparam>LABEL_TEXT no</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>112</ID>
<type>AA_LABEL</type>
<position>53,-50</position>
<gparam>LABEL_TEXT x</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>113</ID>
<type>AA_LABEL</type>
<position>53.5,-83.5</position>
<gparam>LABEL_TEXT y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>114</ID>
<type>GA_LED</type>
<position>137.5,-62.5</position>
<input>
<ID>N_in0</ID>82 </input>
<input>
<ID>N_in1</ID>121 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>118</ID>
<type>AA_LABEL</type>
<position>74.5,-53.5</position>
<gparam>LABEL_TEXT if zx then make x be zero</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>119</ID>
<type>AA_FULLADDER_1BIT</type>
<position>130,-62.5</position>
<input>
<ID>IN_0</ID>120 </input>
<input>
<ID>IN_B_0</ID>119 </input>
<output>
<ID>OUT_0</ID>82 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>120</ID>
<type>AA_LABEL</type>
<position>103.5,-52.5</position>
<gparam>LABEL_TEXT if nx then negate zxo</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>125</ID>
<type>GA_LED</type>
<position>185,-71</position>
<input>
<ID>N_in0</ID>88 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>128</ID>
<type>AA_AND2</type>
<position>131,-79.5</position>
<input>
<ID>IN_0</ID>120 </input>
<input>
<ID>IN_1</ID>119 </input>
<output>
<ID>OUT</ID>83 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>129</ID>
<type>GA_LED</type>
<position>137.5,-79.5</position>
<input>
<ID>N_in0</ID>83 </input>
<input>
<ID>N_in1</ID>122 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>130</ID>
<type>AA_LABEL</type>
<position>130,-57</position>
<gparam>LABEL_TEXT xo plus yo</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>131</ID>
<type>AA_LABEL</type>
<position>133.5,-74.5</position>
<gparam>LABEL_TEXT xo and yo</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>132</ID>
<type>AA_MUX_2x1</type>
<position>148,-72</position>
<input>
<ID>IN_0</ID>122 </input>
<input>
<ID>IN_1</ID>121 </input>
<output>
<ID>OUT</ID>90 </output>
<input>
<ID>SEL_0</ID>86 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>133</ID>
<type>AA_MUX_2x1</type>
<position>170.5,-71</position>
<input>
<ID>IN_0</ID>127 </input>
<input>
<ID>IN_1</ID>126 </input>
<output>
<ID>OUT</ID>88 </output>
<input>
<ID>SEL_0</ID>89 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>135</ID>
<type>GA_LED</type>
<position>153,-72</position>
<input>
<ID>N_in0</ID>90 </input>
<input>
<ID>N_in1</ID>127 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>139</ID>
<type>AA_MUX_2x1</type>
<position>79.5,-48</position>
<input>
<ID>IN_0</ID>100 </input>
<input>
<ID>IN_1</ID>101 </input>
<output>
<ID>OUT</ID>95 </output>
<input>
<ID>SEL_0</ID>99 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>141</ID>
<type>GA_LED</type>
<position>85.5,-48</position>
<input>
<ID>N_in0</ID>95 </input>
<input>
<ID>N_in1</ID>129 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>143</ID>
<type>FF_GND</type>
<position>56.5,-45</position>
<output>
<ID>OUT_0</ID>101 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>151</ID>
<type>AA_MUX_2x1</type>
<position>73.5,-83</position>
<input>
<ID>IN_0</ID>105 </input>
<input>
<ID>IN_1</ID>106 </input>
<output>
<ID>OUT</ID>109 </output>
<input>
<ID>SEL_0</ID>108 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>153</ID>
<type>FF_GND</type>
<position>56,-79.5</position>
<output>
<ID>OUT_0</ID>106 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>155</ID>
<type>GA_LED</type>
<position>79,-83</position>
<input>
<ID>N_in0</ID>109 </input>
<input>
<ID>N_in1</ID>132 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>170</ID>
<type>AA_LABEL</type>
<position>179,-67.5</position>
<gparam>LABEL_TEXT if no then negate fo</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>172</ID>
<type>AA_INVERTER</type>
<position>162,-67</position>
<input>
<ID>IN_0</ID>127 </input>
<output>
<ID>OUT_0</ID>126 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>174</ID>
<type>AA_MUX_2x1</type>
<position>102.5,-47</position>
<input>
<ID>IN_0</ID>129 </input>
<input>
<ID>IN_1</ID>128 </input>
<output>
<ID>OUT</ID>131 </output>
<input>
<ID>SEL_0</ID>130 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>176</ID>
<type>AA_INVERTER</type>
<position>93.5,-44.5</position>
<input>
<ID>IN_0</ID>129 </input>
<output>
<ID>OUT_0</ID>128 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>178</ID>
<type>GA_LED</type>
<position>108,-47</position>
<input>
<ID>N_in0</ID>131 </input>
<input>
<ID>N_in1</ID>120 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>180</ID>
<type>AA_INVERTER</type>
<position>87.5,-80</position>
<input>
<ID>IN_0</ID>132 </input>
<output>
<ID>OUT_0</ID>133 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>182</ID>
<type>AA_MUX_2x1</type>
<position>96,-82</position>
<input>
<ID>IN_0</ID>132 </input>
<input>
<ID>IN_1</ID>133 </input>
<output>
<ID>OUT</ID>135 </output>
<input>
<ID>SEL_0</ID>134 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>184</ID>
<type>GA_LED</type>
<position>101.5,-82</position>
<input>
<ID>N_in0</ID>135 </input>
<input>
<ID>N_in1</ID>119 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>82</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133,-62.5,136.5,-62.5</points>
<connection>
<GID>114</GID>
<name>N_in0</name></connection>
<connection>
<GID>119</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>134,-79.5,136.5,-79.5</points>
<connection>
<GID>128</GID>
<name>OUT</name></connection>
<connection>
<GID>129</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>148,-69.5,148,-28.5</points>
<connection>
<GID>132</GID>
<name>SEL_0</name></connection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>144.5,-28.5,148,-28.5</points>
<connection>
<GID>101</GID>
<name>OUT_0</name></connection>
<intersection>148 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>172.5,-71,184,-71</points>
<connection>
<GID>133</GID>
<name>OUT</name></connection>
<connection>
<GID>125</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170.5,-68.5,170.5,-28.5</points>
<connection>
<GID>133</GID>
<name>SEL_0</name></connection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>158,-28.5,170.5,-28.5</points>
<connection>
<GID>102</GID>
<name>OUT_0</name></connection>
<intersection>170.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>150,-72,152,-72</points>
<connection>
<GID>132</GID>
<name>OUT</name></connection>
<connection>
<GID>135</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>81.5,-48,84.5,-48</points>
<connection>
<GID>139</GID>
<name>OUT</name></connection>
<connection>
<GID>141</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79.5,-45.5,79.5,-30</points>
<connection>
<GID>139</GID>
<name>SEL_0</name></connection>
<intersection>-30 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>71.5,-30,79.5,-30</points>
<connection>
<GID>94</GID>
<name>OUT_0</name></connection>
<intersection>79.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,-51,63.5,-49</points>
<intersection>-51 2</intersection>
<intersection>-49 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>63.5,-49,77.5,-49</points>
<connection>
<GID>139</GID>
<name>IN_0</name></connection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>58.5,-51,63.5,-51</points>
<connection>
<GID>103</GID>
<name>OUT_0</name></connection>
<intersection>63.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68,-47,68,-44</points>
<intersection>-47 1</intersection>
<intersection>-44 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>68,-47,77.5,-47</points>
<connection>
<GID>139</GID>
<name>IN_1</name></connection>
<intersection>68 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56.5,-44,68,-44</points>
<connection>
<GID>143</GID>
<name>OUT_0</name></connection>
<intersection>68 0</intersection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>58.5,-84,71.5,-84</points>
<connection>
<GID>151</GID>
<name>IN_0</name></connection>
<connection>
<GID>105</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>62.5,-82,62.5,-78.5</points>
<intersection>-82 1</intersection>
<intersection>-78.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62.5,-82,71.5,-82</points>
<connection>
<GID>151</GID>
<name>IN_1</name></connection>
<intersection>62.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>56,-78.5,62.5,-78.5</points>
<connection>
<GID>153</GID>
<name>OUT_0</name></connection>
<intersection>62.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,-80.5,73.5,-68.5</points>
<connection>
<GID>151</GID>
<name>SEL_0</name></connection>
<intersection>-68.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>71,-68.5,73.5,-68.5</points>
<connection>
<GID>99</GID>
<name>OUT_0</name></connection>
<intersection>73.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75.5,-83,78,-83</points>
<connection>
<GID>155</GID>
<name>N_in0</name></connection>
<connection>
<GID>151</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>119</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118,-82,118,-63.5</points>
<intersection>-82 5</intersection>
<intersection>-80.5 4</intersection>
<intersection>-63.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>118,-63.5,127,-63.5</points>
<connection>
<GID>119</GID>
<name>IN_B_0</name></connection>
<intersection>118 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>118,-80.5,128,-80.5</points>
<connection>
<GID>128</GID>
<name>IN_1</name></connection>
<intersection>118 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>102.5,-82,118,-82</points>
<connection>
<GID>184</GID>
<name>N_in1</name></connection>
<intersection>118 0</intersection></hsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118,-78.5,118,-47</points>
<intersection>-78.5 3</intersection>
<intersection>-61.5 1</intersection>
<intersection>-47 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>118,-61.5,127,-61.5</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>118 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>118,-78.5,128,-78.5</points>
<connection>
<GID>128</GID>
<name>IN_0</name></connection>
<intersection>118 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>109,-47,118,-47</points>
<connection>
<GID>178</GID>
<name>N_in1</name></connection>
<intersection>118 0</intersection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-71,142,-62.5</points>
<intersection>-71 2</intersection>
<intersection>-62.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138.5,-62.5,142,-62.5</points>
<connection>
<GID>114</GID>
<name>N_in1</name></connection>
<intersection>142 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>142,-71,146,-71</points>
<connection>
<GID>132</GID>
<name>IN_1</name></connection>
<intersection>142 0</intersection></hsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>142,-79.5,142,-73</points>
<intersection>-79.5 1</intersection>
<intersection>-73 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138.5,-79.5,142,-79.5</points>
<connection>
<GID>129</GID>
<name>N_in1</name></connection>
<intersection>142 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>142,-73,146,-73</points>
<connection>
<GID>132</GID>
<name>IN_0</name></connection>
<intersection>142 0</intersection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>167,-70,167,-67</points>
<intersection>-70 2</intersection>
<intersection>-67 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>165,-67,167,-67</points>
<connection>
<GID>172</GID>
<name>OUT_0</name></connection>
<intersection>167 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>167,-70,168.5,-70</points>
<connection>
<GID>133</GID>
<name>IN_1</name></connection>
<intersection>167 0</intersection></hsegment></shape></wire>
<wire>
<ID>127</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156.5,-72,156.5,-67</points>
<intersection>-72 2</intersection>
<intersection>-67 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>156.5,-67,159,-67</points>
<connection>
<GID>172</GID>
<name>IN_0</name></connection>
<intersection>156.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>154,-72,168.5,-72</points>
<connection>
<GID>135</GID>
<name>N_in1</name></connection>
<connection>
<GID>133</GID>
<name>IN_0</name></connection>
<intersection>156.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>128</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97.5,-46,97.5,-44.5</points>
<intersection>-46 2</intersection>
<intersection>-44.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>96.5,-44.5,97.5,-44.5</points>
<connection>
<GID>176</GID>
<name>OUT_0</name></connection>
<intersection>97.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97.5,-46,100.5,-46</points>
<connection>
<GID>174</GID>
<name>IN_1</name></connection>
<intersection>97.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>129</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>86.5,-48,100.5,-48</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<connection>
<GID>141</GID>
<name>N_in1</name></connection>
<intersection>90.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>90.5,-48,90.5,-44.5</points>
<connection>
<GID>176</GID>
<name>IN_0</name></connection>
<intersection>-48 1</intersection></vsegment></shape></wire>
<wire>
<ID>130</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102.5,-44.5,102.5,-30</points>
<connection>
<GID>174</GID>
<name>SEL_0</name></connection>
<intersection>-30 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>90.5,-30,102.5,-30</points>
<connection>
<GID>96</GID>
<name>OUT_0</name></connection>
<intersection>102.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104.5,-47,107,-47</points>
<connection>
<GID>178</GID>
<name>N_in0</name></connection>
<connection>
<GID>174</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>80,-83,94,-83</points>
<connection>
<GID>155</GID>
<name>N_in1</name></connection>
<connection>
<GID>182</GID>
<name>IN_0</name></connection>
<intersection>84.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>84.5,-83,84.5,-80</points>
<connection>
<GID>180</GID>
<name>IN_0</name></connection>
<intersection>-83 1</intersection></vsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>92,-81,92,-80</points>
<intersection>-81 1</intersection>
<intersection>-80 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>92,-81,94,-81</points>
<connection>
<GID>182</GID>
<name>IN_1</name></connection>
<intersection>92 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-80,92,-80</points>
<connection>
<GID>180</GID>
<name>OUT_0</name></connection>
<intersection>92 0</intersection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96,-79.5,96,-68.5</points>
<connection>
<GID>182</GID>
<name>SEL_0</name></connection>
<intersection>-68.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85.5,-68.5,96,-68.5</points>
<connection>
<GID>100</GID>
<name>OUT_0</name></connection>
<intersection>96 0</intersection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>98,-82,100.5,-82</points>
<connection>
<GID>184</GID>
<name>N_in0</name></connection>
<connection>
<GID>182</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>172.568,-23.7705,295.958,-85.9082</PageViewport>
<gate>
<ID>193</ID>
<type>AA_TOGGLE</type>
<position>93.5,-32.5</position>
<output>
<ID>OUT_0</ID>144 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>194</ID>
<type>AA_LABEL</type>
<position>189.5,-57.5</position>
<gparam>LABEL_TEXT if f then xo+yo else xo&yo</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>195</ID>
<type>AA_TOGGLE</type>
<position>93.5,-65.5</position>
<output>
<ID>OUT_0</ID>146 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>3</ID>
<type>AE_OR2</type>
<position>229,-59</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>196</ID>
<type>AA_LABEL</type>
<position>107,-7.5</position>
<gparam>LABEL_TEXT zx</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>197</ID>
<type>AA_LABEL</type>
<position>126,-7.5</position>
<gparam>LABEL_TEXT nx</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>198</ID>
<type>AA_LABEL</type>
<position>106.5,-46</position>
<gparam>LABEL_TEXT zy</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>199</ID>
<type>AA_LABEL</type>
<position>121,-46</position>
<gparam>LABEL_TEXT ny</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>200</ID>
<type>AA_LABEL</type>
<position>179.5,-6</position>
<gparam>LABEL_TEXT f</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>201</ID>
<type>AA_LABEL</type>
<position>193,-6.5</position>
<gparam>LABEL_TEXT no</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>202</ID>
<type>AA_LABEL</type>
<position>90,-31.5</position>
<gparam>LABEL_TEXT x</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>203</ID>
<type>AA_LABEL</type>
<position>90.5,-65</position>
<gparam>LABEL_TEXT y</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>204</ID>
<type>GA_LED</type>
<position>174.5,-44</position>
<input>
<ID>N_in0</ID>136 </input>
<input>
<ID>N_in1</ID>152 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>205</ID>
<type>AA_LABEL</type>
<position>111.5,-35</position>
<gparam>LABEL_TEXT if zx then make x be zero</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>206</ID>
<type>AA_FULLADDER_1BIT</type>
<position>167,-44</position>
<input>
<ID>IN_0</ID>151 </input>
<input>
<ID>IN_B_0</ID>150 </input>
<output>
<ID>OUT_0</ID>136 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>207</ID>
<type>AA_LABEL</type>
<position>140.5,-34</position>
<gparam>LABEL_TEXT if nx then negate zxo</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>208</ID>
<type>GA_LED</type>
<position>216,-52.5</position>
<input>
<ID>N_in0</ID>139 </input>
<input>
<ID>N_in1</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>209</ID>
<type>AA_AND2</type>
<position>168,-61</position>
<input>
<ID>IN_0</ID>151 </input>
<input>
<ID>IN_1</ID>150 </input>
<output>
<ID>OUT</ID>137 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>210</ID>
<type>GA_LED</type>
<position>174.5,-61</position>
<input>
<ID>N_in0</ID>137 </input>
<input>
<ID>N_in1</ID>153 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>211</ID>
<type>AA_LABEL</type>
<position>167,-38.5</position>
<gparam>LABEL_TEXT xo plus yo</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>212</ID>
<type>AA_LABEL</type>
<position>170.5,-56</position>
<gparam>LABEL_TEXT xo and yo</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>213</ID>
<type>AA_MUX_2x1</type>
<position>185,-53.5</position>
<input>
<ID>IN_0</ID>153 </input>
<input>
<ID>IN_1</ID>152 </input>
<output>
<ID>OUT</ID>141 </output>
<input>
<ID>SEL_0</ID>138 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>21</ID>
<type>AA_INVERTER</type>
<position>238,-59</position>
<input>
<ID>IN_0</ID>7 </input>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>214</ID>
<type>AA_MUX_2x1</type>
<position>207.5,-52.5</position>
<input>
<ID>IN_0</ID>155 </input>
<input>
<ID>IN_1</ID>154 </input>
<output>
<ID>OUT</ID>139 </output>
<input>
<ID>SEL_0</ID>140 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>215</ID>
<type>GA_LED</type>
<position>190,-53.5</position>
<input>
<ID>N_in0</ID>141 </input>
<input>
<ID>N_in1</ID>155 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>216</ID>
<type>AA_MUX_2x1</type>
<position>116.5,-29.5</position>
<input>
<ID>IN_0</ID>144 </input>
<input>
<ID>IN_1</ID>145 </input>
<output>
<ID>OUT</ID>142 </output>
<input>
<ID>SEL_0</ID>143 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>217</ID>
<type>GA_LED</type>
<position>122.5,-29.5</position>
<input>
<ID>N_in0</ID>142 </input>
<input>
<ID>N_in1</ID>157 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>218</ID>
<type>FF_GND</type>
<position>93.5,-26.5</position>
<output>
<ID>OUT_0</ID>145 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>219</ID>
<type>AA_MUX_2x1</type>
<position>110.5,-64.5</position>
<input>
<ID>IN_0</ID>146 </input>
<input>
<ID>IN_1</ID>147 </input>
<output>
<ID>OUT</ID>149 </output>
<input>
<ID>SEL_0</ID>148 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>27</ID>
<type>GA_LED</type>
<position>243.5,-59</position>
<input>
<ID>N_in0</ID>13 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>220</ID>
<type>FF_GND</type>
<position>93,-61</position>
<output>
<ID>OUT_0</ID>147 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>221</ID>
<type>GA_LED</type>
<position>116,-64.5</position>
<input>
<ID>N_in0</ID>149 </input>
<input>
<ID>N_in1</ID>160 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>222</ID>
<type>AA_LABEL</type>
<position>216,-49</position>
<gparam>LABEL_TEXT if no then negate fo</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>223</ID>
<type>AA_INVERTER</type>
<position>199,-48.5</position>
<input>
<ID>IN_0</ID>155 </input>
<output>
<ID>OUT_0</ID>154 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>224</ID>
<type>AA_MUX_2x1</type>
<position>139.5,-28.5</position>
<input>
<ID>IN_0</ID>157 </input>
<input>
<ID>IN_1</ID>156 </input>
<output>
<ID>OUT</ID>159 </output>
<input>
<ID>SEL_0</ID>158 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>225</ID>
<type>AA_INVERTER</type>
<position>130.5,-26</position>
<input>
<ID>IN_0</ID>157 </input>
<output>
<ID>OUT_0</ID>156 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>226</ID>
<type>GA_LED</type>
<position>145,-28.5</position>
<input>
<ID>N_in0</ID>159 </input>
<input>
<ID>N_in1</ID>151 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>227</ID>
<type>AA_INVERTER</type>
<position>124.5,-61.5</position>
<input>
<ID>IN_0</ID>160 </input>
<output>
<ID>OUT_0</ID>161 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>228</ID>
<type>AA_MUX_2x1</type>
<position>133,-63.5</position>
<input>
<ID>IN_0</ID>160 </input>
<input>
<ID>IN_1</ID>161 </input>
<output>
<ID>OUT</ID>163 </output>
<input>
<ID>SEL_0</ID>162 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>229</ID>
<type>GA_LED</type>
<position>138.5,-63.5</position>
<input>
<ID>N_in0</ID>163 </input>
<input>
<ID>N_in1</ID>150 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>231</ID>
<type>AA_LABEL</type>
<position>234,-64</position>
<gparam>LABEL_TEXT if out=0 then zr = 1 else zr = 0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>233</ID>
<type>FF_GND</type>
<position>219.5,-69</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>185</ID>
<type>AA_LABEL</type>
<position>106,-69.5</position>
<gparam>LABEL_TEXT if zy then make y be zero</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>186</ID>
<type>AA_LABEL</type>
<position>133.5,-69</position>
<gparam>LABEL_TEXT if ny then negate zyo</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>187</ID>
<type>AA_TOGGLE</type>
<position>106.5,-11.5</position>
<output>
<ID>OUT_0</ID>143 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>188</ID>
<type>AA_TOGGLE</type>
<position>125.5,-11.5</position>
<output>
<ID>OUT_0</ID>158 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>189</ID>
<type>AA_TOGGLE</type>
<position>106,-50</position>
<output>
<ID>OUT_0</ID>148 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>190</ID>
<type>AA_TOGGLE</type>
<position>120.5,-50</position>
<output>
<ID>OUT_0</ID>162 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>191</ID>
<type>AA_TOGGLE</type>
<position>179.5,-10</position>
<output>
<ID>OUT_0</ID>138 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>192</ID>
<type>AA_TOGGLE</type>
<position>193,-10</position>
<output>
<ID>OUT_0</ID>140 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>219.5,-58,226,-58</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>219.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>219.5,-58,219.5,-52.5</points>
<intersection>-58 1</intersection>
<intersection>-52.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>217,-52.5,219.5,-52.5</points>
<connection>
<GID>208</GID>
<name>N_in1</name></connection>
<intersection>219.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>232,-59,235,-59</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<connection>
<GID>3</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>241,-59,242.5,-59</points>
<connection>
<GID>27</GID>
<name>N_in0</name></connection>
<connection>
<GID>21</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>219.5,-68,219.5,-60</points>
<connection>
<GID>233</GID>
<name>OUT_0</name></connection>
<intersection>-60 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>219.5,-60,226,-60</points>
<connection>
<GID>3</GID>
<name>IN_1</name></connection>
<intersection>219.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>170,-44,173.5,-44</points>
<connection>
<GID>206</GID>
<name>OUT_0</name></connection>
<connection>
<GID>204</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>171,-61,173.5,-61</points>
<connection>
<GID>209</GID>
<name>OUT</name></connection>
<connection>
<GID>210</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>185,-51,185,-10</points>
<connection>
<GID>213</GID>
<name>SEL_0</name></connection>
<intersection>-10 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>181.5,-10,185,-10</points>
<connection>
<GID>191</GID>
<name>OUT_0</name></connection>
<intersection>185 0</intersection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>209.5,-52.5,215,-52.5</points>
<connection>
<GID>214</GID>
<name>OUT</name></connection>
<connection>
<GID>208</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>140</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207.5,-50,207.5,-10</points>
<connection>
<GID>214</GID>
<name>SEL_0</name></connection>
<intersection>-10 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>195,-10,207.5,-10</points>
<connection>
<GID>192</GID>
<name>OUT_0</name></connection>
<intersection>207.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<hsegment>
<ID>5</ID>
<points>187,-53.5,189,-53.5</points>
<connection>
<GID>213</GID>
<name>OUT</name></connection>
<connection>
<GID>215</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>142</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>118.5,-29.5,121.5,-29.5</points>
<connection>
<GID>216</GID>
<name>OUT</name></connection>
<connection>
<GID>217</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>143</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,-27,116.5,-11.5</points>
<connection>
<GID>216</GID>
<name>SEL_0</name></connection>
<intersection>-11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108.5,-11.5,116.5,-11.5</points>
<connection>
<GID>187</GID>
<name>OUT_0</name></connection>
<intersection>116.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>144</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100.5,-32.5,100.5,-30.5</points>
<intersection>-32.5 2</intersection>
<intersection>-30.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>100.5,-30.5,114.5,-30.5</points>
<connection>
<GID>216</GID>
<name>IN_0</name></connection>
<intersection>100.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>95.5,-32.5,100.5,-32.5</points>
<connection>
<GID>193</GID>
<name>OUT_0</name></connection>
<intersection>100.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>145</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>105,-28.5,105,-25.5</points>
<intersection>-28.5 1</intersection>
<intersection>-25.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>105,-28.5,114.5,-28.5</points>
<connection>
<GID>216</GID>
<name>IN_1</name></connection>
<intersection>105 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>93.5,-25.5,105,-25.5</points>
<connection>
<GID>218</GID>
<name>OUT_0</name></connection>
<intersection>105 0</intersection></hsegment></shape></wire>
<wire>
<ID>146</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>95.5,-65.5,108.5,-65.5</points>
<connection>
<GID>195</GID>
<name>OUT_0</name></connection>
<connection>
<GID>219</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>147</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99.5,-63.5,99.5,-60</points>
<intersection>-63.5 1</intersection>
<intersection>-60 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>99.5,-63.5,108.5,-63.5</points>
<connection>
<GID>219</GID>
<name>IN_1</name></connection>
<intersection>99.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>93,-60,99.5,-60</points>
<connection>
<GID>220</GID>
<name>OUT_0</name></connection>
<intersection>99.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>148</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>110.5,-62,110.5,-50</points>
<connection>
<GID>219</GID>
<name>SEL_0</name></connection>
<intersection>-50 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>108,-50,110.5,-50</points>
<connection>
<GID>189</GID>
<name>OUT_0</name></connection>
<intersection>110.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>149</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>112.5,-64.5,115,-64.5</points>
<connection>
<GID>219</GID>
<name>OUT</name></connection>
<connection>
<GID>221</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>150</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155,-63.5,155,-45</points>
<intersection>-63.5 5</intersection>
<intersection>-62 4</intersection>
<intersection>-45 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>155,-45,164,-45</points>
<connection>
<GID>206</GID>
<name>IN_B_0</name></connection>
<intersection>155 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>155,-62,165,-62</points>
<connection>
<GID>209</GID>
<name>IN_1</name></connection>
<intersection>155 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>139.5,-63.5,155,-63.5</points>
<connection>
<GID>229</GID>
<name>N_in1</name></connection>
<intersection>155 0</intersection></hsegment></shape></wire>
<wire>
<ID>151</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>155,-60,155,-28.5</points>
<intersection>-60 3</intersection>
<intersection>-43 1</intersection>
<intersection>-28.5 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>155,-43,164,-43</points>
<connection>
<GID>206</GID>
<name>IN_0</name></connection>
<intersection>155 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>155,-60,165,-60</points>
<connection>
<GID>209</GID>
<name>IN_0</name></connection>
<intersection>155 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>146,-28.5,155,-28.5</points>
<connection>
<GID>226</GID>
<name>N_in1</name></connection>
<intersection>155 0</intersection></hsegment></shape></wire>
<wire>
<ID>152</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179,-52.5,179,-44</points>
<intersection>-52.5 2</intersection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>175.5,-44,179,-44</points>
<connection>
<GID>204</GID>
<name>N_in1</name></connection>
<intersection>179 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>179,-52.5,183,-52.5</points>
<connection>
<GID>213</GID>
<name>IN_1</name></connection>
<intersection>179 0</intersection></hsegment></shape></wire>
<wire>
<ID>153</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>179,-61,179,-54.5</points>
<intersection>-61 1</intersection>
<intersection>-54.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>175.5,-61,179,-61</points>
<connection>
<GID>210</GID>
<name>N_in1</name></connection>
<intersection>179 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>179,-54.5,183,-54.5</points>
<connection>
<GID>213</GID>
<name>IN_0</name></connection>
<intersection>179 0</intersection></hsegment></shape></wire>
<wire>
<ID>154</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>204,-51.5,204,-48.5</points>
<intersection>-51.5 2</intersection>
<intersection>-48.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>202,-48.5,204,-48.5</points>
<connection>
<GID>223</GID>
<name>OUT_0</name></connection>
<intersection>204 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>204,-51.5,205.5,-51.5</points>
<connection>
<GID>214</GID>
<name>IN_1</name></connection>
<intersection>204 0</intersection></hsegment></shape></wire>
<wire>
<ID>155</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>193.5,-53.5,193.5,-48.5</points>
<intersection>-53.5 2</intersection>
<intersection>-48.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>193.5,-48.5,196,-48.5</points>
<connection>
<GID>223</GID>
<name>IN_0</name></connection>
<intersection>193.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>191,-53.5,205.5,-53.5</points>
<connection>
<GID>214</GID>
<name>IN_0</name></connection>
<connection>
<GID>215</GID>
<name>N_in1</name></connection>
<intersection>193.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>156</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>134.5,-27.5,134.5,-26</points>
<intersection>-27.5 2</intersection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>133.5,-26,134.5,-26</points>
<connection>
<GID>225</GID>
<name>OUT_0</name></connection>
<intersection>134.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>134.5,-27.5,137.5,-27.5</points>
<connection>
<GID>224</GID>
<name>IN_1</name></connection>
<intersection>134.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>157</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>123.5,-29.5,137.5,-29.5</points>
<connection>
<GID>217</GID>
<name>N_in1</name></connection>
<connection>
<GID>224</GID>
<name>IN_0</name></connection>
<intersection>127.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>127.5,-29.5,127.5,-26</points>
<connection>
<GID>225</GID>
<name>IN_0</name></connection>
<intersection>-29.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>158</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>139.5,-26,139.5,-11.5</points>
<connection>
<GID>224</GID>
<name>SEL_0</name></connection>
<intersection>-11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>127.5,-11.5,139.5,-11.5</points>
<connection>
<GID>188</GID>
<name>OUT_0</name></connection>
<intersection>139.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>159</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>141.5,-28.5,144,-28.5</points>
<connection>
<GID>224</GID>
<name>OUT</name></connection>
<connection>
<GID>226</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>160</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>117,-64.5,131,-64.5</points>
<connection>
<GID>221</GID>
<name>N_in1</name></connection>
<connection>
<GID>228</GID>
<name>IN_0</name></connection>
<intersection>121.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>121.5,-64.5,121.5,-61.5</points>
<connection>
<GID>227</GID>
<name>IN_0</name></connection>
<intersection>-64.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>161</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129,-62.5,129,-61.5</points>
<intersection>-62.5 1</intersection>
<intersection>-61.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>129,-62.5,131,-62.5</points>
<connection>
<GID>228</GID>
<name>IN_1</name></connection>
<intersection>129 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>127.5,-61.5,129,-61.5</points>
<connection>
<GID>227</GID>
<name>OUT_0</name></connection>
<intersection>129 0</intersection></hsegment></shape></wire>
<wire>
<ID>162</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,-61,133,-50</points>
<connection>
<GID>228</GID>
<name>SEL_0</name></connection>
<intersection>-50 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>122.5,-50,133,-50</points>
<connection>
<GID>190</GID>
<name>OUT_0</name></connection>
<intersection>133 0</intersection></hsegment></shape></wire>
<wire>
<ID>163</ID>
<shape>
<hsegment>
<ID>3</ID>
<points>135,-63.5,137.5,-63.5</points>
<connection>
<GID>228</GID>
<name>OUT</name></connection>
<connection>
<GID>229</GID>
<name>N_in0</name></connection></hsegment></shape></wire></page 2>
<page 3>
<PageViewport>-5.90755,60.8509,323.133,-104.85</PageViewport>
<gate>
<ID>249</ID>
<type>AA_TOGGLE</type>
<position>22.5,11</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>251</ID>
<type>AA_TOGGLE</type>
<position>22.5,8</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>253</ID>
<type>AA_TOGGLE</type>
<position>22,5</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>255</ID>
<type>AA_TOGGLE</type>
<position>22.5,2</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>257</ID>
<type>AA_LABEL</type>
<position>24,15</position>
<gparam>LABEL_TEXT A bus</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>258</ID>
<type>AA_TOGGLE</type>
<position>22,-5.5</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>259</ID>
<type>AA_TOGGLE</type>
<position>22,-8.5</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>260</ID>
<type>AA_TOGGLE</type>
<position>21.5,-11.5</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>261</ID>
<type>AA_TOGGLE</type>
<position>22,-14.5</position>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>262</ID>
<type>AA_LABEL</type>
<position>23.5,-1.5</position>
<gparam>LABEL_TEXT B bus</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>264</ID>
<type>AA_LABEL</type>
<position>17.5,11.5</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>265</ID>
<type>AA_LABEL</type>
<position>17.5,8</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>266</ID>
<type>AA_LABEL</type>
<position>17.5,5</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>267</ID>
<type>AA_LABEL</type>
<position>17.5,2</position>
<gparam>LABEL_TEXT 3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>268</ID>
<type>AA_LABEL</type>
<position>17.5,-5</position>
<gparam>LABEL_TEXT 0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>269</ID>
<type>AA_LABEL</type>
<position>17.5,-8.5</position>
<gparam>LABEL_TEXT 1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>270</ID>
<type>AA_LABEL</type>
<position>17.5,-11.5</position>
<gparam>LABEL_TEXT 2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>271</ID>
<type>AA_LABEL</type>
<position>17.5,-14.5</position>
<gparam>LABEL_TEXT 3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>272</ID>
<type>AA_LABEL</type>
<position>23.5,24.5</position>
<gparam>LABEL_TEXT out</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate></page 3>
<page 4>
<PageViewport>0,156.824,1386.58,-541.438</PageViewport></page 4>
<page 5>
<PageViewport>0,156.824,1386.58,-541.438</PageViewport></page 5>
<page 6>
<PageViewport>0,156.824,1386.58,-541.438</PageViewport></page 6>
<page 7>
<PageViewport>0,156.824,1386.58,-541.438</PageViewport></page 7>
<page 8>
<PageViewport>0,156.824,1386.58,-541.438</PageViewport></page 8>
<page 9>
<PageViewport>0,156.824,1386.58,-541.438</PageViewport></page 9></circuit>